magic
tech sky130A
magscale 1 2
timestamp 1770389962
<< viali >>
rect 4362 -990 4810 -906
rect 8348 -974 8798 -906
rect 12304 -1002 12744 -924
rect 68398 -10766 68446 -10620
rect 74044 -10758 74146 -10622
rect 60058 -11876 60094 -11754
rect 64180 -11922 64244 -11796
rect 70034 -11940 70090 -11808
rect 73440 -11948 73496 -11816
rect 4116 -22706 4522 -22660
rect 8296 -22706 8646 -22644
rect 12778 -22738 13126 -22670
<< metal1 >>
rect 15604 15128 31505 15902
rect 46628 15058 63915 15832
rect -266 9686 126 9822
rect -276 9474 126 9686
rect -266 9300 126 9474
rect -2524 6645 -1875 6649
rect -952 6645 344 6722
rect -2524 6466 344 6645
rect -2524 -4323 -2345 6466
rect -952 6454 344 6466
rect -952 6278 -704 6454
rect -952 6238 -703 6278
rect -941 -981 -703 6238
rect 4358 -900 4814 178
rect 8350 -900 8802 128
rect 4350 -906 4822 -900
rect -941 -1010 1493 -981
rect 4350 -990 4362 -906
rect 4810 -990 4822 -906
rect 8336 -906 8810 -900
rect 8336 -974 8348 -906
rect 8798 -974 8810 -906
rect 12308 -918 12750 82
rect 15153 4 31629 766
rect 46628 -66 63671 696
rect 8336 -980 8810 -974
rect 12292 -924 12756 -918
rect 8350 -982 8802 -980
rect 4350 -996 4822 -990
rect -941 -1216 3290 -1010
rect 5758 -1182 7214 -1008
rect 9810 -1190 11334 -996
rect 12292 -1002 12304 -924
rect 12744 -1002 12756 -924
rect 12292 -1008 12756 -1002
rect 13838 -1182 15690 -1016
rect -941 -1219 1493 -1216
rect -2518 -4560 -2352 -4323
rect -3788 -5620 -3411 -5618
rect -2518 -5620 -2356 -5064
rect -3788 -5776 -2356 -5620
rect -3790 -5804 -2356 -5776
rect -3790 -5884 -3410 -5804
rect -3790 -6058 -3404 -5884
rect -3790 -6680 -3410 -6058
rect -2518 -6372 -2356 -5804
rect -3782 -33342 -3415 -6680
rect -2554 -15577 -2375 -6786
rect 15337 -7058 31489 -6284
rect 74241 -10604 74432 -10602
rect 68410 -10608 69882 -10604
rect 68392 -10620 69882 -10608
rect 57939 -11095 58237 -10653
rect 56580 -11393 58237 -11095
rect 64123 -11105 64421 -10657
rect 56580 -11848 56878 -11393
rect 62734 -11403 64421 -11105
rect 66546 -11149 66844 -11139
rect 67947 -11149 68245 -10671
rect 68392 -10766 68398 -10620
rect 68446 -10766 69882 -10620
rect 74038 -10612 74152 -10610
rect 74202 -10612 74432 -10604
rect 74038 -10622 74432 -10612
rect 68392 -10778 69882 -10766
rect 68410 -10784 69882 -10778
rect 60052 -11750 60100 -11742
rect 59642 -11754 60210 -11750
rect 59642 -11876 60058 -11754
rect 60094 -11876 60210 -11754
rect 62734 -11858 63032 -11403
rect 66546 -11447 68245 -11149
rect 64174 -11792 64250 -11784
rect 63780 -11796 64328 -11792
rect 59642 -13147 60210 -11876
rect 63780 -11922 64180 -11796
rect 64244 -11922 64328 -11796
rect 66546 -11892 66844 -11447
rect 69704 -11798 69881 -10784
rect 73597 -11135 73895 -10683
rect 74038 -10758 74044 -10622
rect 74146 -10758 74432 -10622
rect 74038 -10770 74432 -10758
rect 74082 -10772 74432 -10770
rect 74202 -10808 74432 -10772
rect 72276 -11433 73895 -11135
rect 70028 -11798 70096 -11796
rect 69608 -11808 70116 -11798
rect 63780 -13147 64328 -11922
rect 69608 -11940 70034 -11808
rect 70090 -11940 70116 -11808
rect 72276 -11892 72574 -11433
rect 73434 -11816 73502 -11804
rect 73434 -11818 73440 -11816
rect 69608 -13147 70116 -11940
rect 73024 -11948 73440 -11818
rect 73496 -11948 73502 -11816
rect 73024 -11960 73502 -11948
rect 73024 -13147 73470 -11960
rect 74241 -13147 74432 -10808
rect 78655 -13147 79417 781
rect 59373 -13909 79417 -13147
rect -960 -15472 18 -15432
rect -960 -15577 292 -15472
rect -2554 -15756 292 -15577
rect -962 -15757 292 -15756
rect -960 -15832 292 -15757
rect -960 -22568 -722 -15832
rect -694 -15834 292 -15832
rect -962 -22706 -716 -22568
rect 4124 -22654 4514 -22092
rect 8302 -22638 8654 -22070
rect 8284 -22644 8658 -22638
rect 4104 -22660 4534 -22654
rect 4104 -22706 4116 -22660
rect 4522 -22706 4534 -22660
rect -976 -22932 2948 -22706
rect 4104 -22712 4534 -22706
rect 8284 -22706 8296 -22644
rect 8646 -22706 8658 -22644
rect 12774 -22664 13134 -22008
rect 15411 -22182 31889 -21420
rect 59373 -21494 60135 -13909
rect 46309 -22256 60135 -21494
rect 8284 -22712 8658 -22706
rect 12766 -22670 13138 -22664
rect 5546 -22922 7314 -22720
rect 12766 -22738 12778 -22670
rect 13126 -22738 13138 -22670
rect 9754 -22940 11832 -22738
rect 12766 -22744 13138 -22738
rect 15169 -28034 31487 -27260
rect -3782 -33657 204 -33342
rect -3774 -33864 204 -33657
rect 15411 -43158 31457 -42396
rect 78655 -42400 79417 -13909
rect 46099 -43162 79417 -42400
use sky130_fd_pr__cap_mim_m3_1_L6ZKLG  sky130_fd_pr__cap_mim_m3_1_L6ZKLG_0
timestamp 1770389351
transform 1 0 70092 0 1 -31238
box -6492 -9480 6492 9480
use OFCB  x1
timestamp 1768581666
transform 1 0 958 0 1 -18688
box -914 -3502 15456 12442
use OFCB  x2
timestamp 1768581666
transform 1 0 31946 0 1 3428
box -914 -3502 15456 12442
use OFCB  x3
timestamp 1768581666
transform 1 0 31844 0 1 -18762
box -914 -3502 15456 12442
use OFCB  x4
timestamp 1768581666
transform 1 0 64098 0 1 3470
box -914 -3502 15456 12442
use OFCB  x5
timestamp 1768581666
transform 1 0 808 0 1 -39664
box -914 -3502 15456 12442
use OFCB  x6
timestamp 1768581666
transform 1 0 31770 0 1 -39668
box -914 -3502 15456 12442
use OFCB  x16
timestamp 1768581666
transform 1 0 922 0 1 3498
box -914 -3502 15456 12442
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR1
timestamp 1770379997
transform 0 1 8508 -1 0 -1089
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR2
timestamp 1770379997
transform 0 1 4324 -1 0 -22827
box -201 -1682 201 1682
use sky130_fd_pr__res_high_po_0p35_NL498X  XR3
timestamp 1770379997
transform 1 0 -2443 0 1 -6616
box -201 -642 201 642
use sky130_fd_pr__res_high_po_0p35_NL498X  XR15
timestamp 1770379997
transform 1 0 -2441 0 1 -4862
box -201 -642 201 642
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR17
timestamp 1770379997
transform 0 1 12576 -1 0 -1107
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR18
timestamp 1770379997
transform 0 1 4552 -1 0 -1107
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR21
timestamp 1770379997
transform 0 1 12936 -1 0 -22847
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR24
timestamp 1770379997
transform 0 1 8496 -1 0 -22827
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR35
timestamp 1770379997
transform 0 1 57384 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR36 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 58230 -1 0 -11817
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR37
timestamp 1770379997
transform 0 1 63554 -1 0 -10683
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_DBPYMX  XR38 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 63371 -1 0 -11857
box -201 -889 201 889
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR39
timestamp 1770379997
transform 0 1 67388 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR40
timestamp 1770379997
transform 0 1 68206 -1 0 -11871
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR41
timestamp 1770379997
transform 0 1 73036 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_MAXMKG  XR42 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 72768 -1 0 -11883
box -201 -742 201 742
<< end >>
