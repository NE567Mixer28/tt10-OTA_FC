magic
tech sky130A
magscale 1 2
timestamp 1770370757
<< metal3 >>
rect -19716 3012 -13344 3040
rect -19716 -3012 -13428 3012
rect -13364 -3012 -13344 3012
rect -19716 -3040 -13344 -3012
rect -13104 3012 -6732 3040
rect -13104 -3012 -6816 3012
rect -6752 -3012 -6732 3012
rect -13104 -3040 -6732 -3012
rect -6492 3012 -120 3040
rect -6492 -3012 -204 3012
rect -140 -3012 -120 3012
rect -6492 -3040 -120 -3012
rect 120 3012 6492 3040
rect 120 -3012 6408 3012
rect 6472 -3012 6492 3012
rect 120 -3040 6492 -3012
rect 6732 3012 13104 3040
rect 6732 -3012 13020 3012
rect 13084 -3012 13104 3012
rect 6732 -3040 13104 -3012
rect 13344 3012 19716 3040
rect 13344 -3012 19632 3012
rect 19696 -3012 19716 3012
rect 13344 -3040 19716 -3012
<< via3 >>
rect -13428 -3012 -13364 3012
rect -6816 -3012 -6752 3012
rect -204 -3012 -140 3012
rect 6408 -3012 6472 3012
rect 13020 -3012 13084 3012
rect 19632 -3012 19696 3012
<< mimcap >>
rect -19676 2960 -13676 3000
rect -19676 -2960 -19636 2960
rect -13716 -2960 -13676 2960
rect -19676 -3000 -13676 -2960
rect -13064 2960 -7064 3000
rect -13064 -2960 -13024 2960
rect -7104 -2960 -7064 2960
rect -13064 -3000 -7064 -2960
rect -6452 2960 -452 3000
rect -6452 -2960 -6412 2960
rect -492 -2960 -452 2960
rect -6452 -3000 -452 -2960
rect 160 2960 6160 3000
rect 160 -2960 200 2960
rect 6120 -2960 6160 2960
rect 160 -3000 6160 -2960
rect 6772 2960 12772 3000
rect 6772 -2960 6812 2960
rect 12732 -2960 12772 2960
rect 6772 -3000 12772 -2960
rect 13384 2960 19384 3000
rect 13384 -2960 13424 2960
rect 19344 -2960 19384 2960
rect 13384 -3000 19384 -2960
<< mimcapcontact >>
rect -19636 -2960 -13716 2960
rect -13024 -2960 -7104 2960
rect -6412 -2960 -492 2960
rect 200 -2960 6120 2960
rect 6812 -2960 12732 2960
rect 13424 -2960 19344 2960
<< metal4 >>
rect -13444 3012 -13348 3028
rect -19637 2960 -13715 2961
rect -19637 -2960 -19636 2960
rect -13716 -2960 -13715 2960
rect -19637 -2961 -13715 -2960
rect -13444 -3012 -13428 3012
rect -13364 -3012 -13348 3012
rect -6832 3012 -6736 3028
rect -13025 2960 -7103 2961
rect -13025 -2960 -13024 2960
rect -7104 -2960 -7103 2960
rect -13025 -2961 -7103 -2960
rect -13444 -3028 -13348 -3012
rect -6832 -3012 -6816 3012
rect -6752 -3012 -6736 3012
rect -220 3012 -124 3028
rect -6413 2960 -491 2961
rect -6413 -2960 -6412 2960
rect -492 -2960 -491 2960
rect -6413 -2961 -491 -2960
rect -6832 -3028 -6736 -3012
rect -220 -3012 -204 3012
rect -140 -3012 -124 3012
rect 6392 3012 6488 3028
rect 199 2960 6121 2961
rect 199 -2960 200 2960
rect 6120 -2960 6121 2960
rect 199 -2961 6121 -2960
rect -220 -3028 -124 -3012
rect 6392 -3012 6408 3012
rect 6472 -3012 6488 3012
rect 13004 3012 13100 3028
rect 6811 2960 12733 2961
rect 6811 -2960 6812 2960
rect 12732 -2960 12733 2960
rect 6811 -2961 12733 -2960
rect 6392 -3028 6488 -3012
rect 13004 -3012 13020 3012
rect 13084 -3012 13100 3012
rect 19616 3012 19712 3028
rect 13423 2960 19345 2961
rect 13423 -2960 13424 2960
rect 19344 -2960 19345 2960
rect 13423 -2961 19345 -2960
rect 13004 -3028 13100 -3012
rect 19616 -3012 19632 3012
rect 19696 -3012 19712 3012
rect 19616 -3028 19712 -3012
<< properties >>
string FIXED_BBOX 13344 -3040 19424 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
