magic
tech sky130A
magscale 1 2
timestamp 1752662732
<< metal1 >>
rect -342 9256 -142 9456
rect 5488 8430 11412 8998
rect 17552 8994 19296 9004
rect 13444 8976 19296 8994
rect 13444 8960 19324 8976
rect 13398 8448 19324 8960
rect 5532 8072 7262 8430
rect 8266 8090 9996 8430
rect 3044 7438 5088 7448
rect 3034 6528 5088 7438
rect -358 5854 -158 6054
rect 3034 5544 3872 6528
rect 7682 6080 7818 8050
rect 6066 5984 6076 6080
rect 6770 5984 6780 6080
rect 8770 5984 8780 6080
rect 9474 5984 9484 6080
rect 3030 4624 5074 5544
rect 3034 4618 3872 4624
rect 7686 4018 7818 5978
rect 10862 4358 11394 8430
rect 13398 8052 15128 8448
rect 16138 8430 19324 8448
rect 16138 8072 17868 8430
rect 13920 5954 13930 6050
rect 14624 5954 14634 6050
rect 16616 5960 16626 6056
rect 17320 5960 17330 6056
rect 6536 3556 7410 3992
rect 9376 3564 10206 3974
rect 10862 3564 11384 4358
rect 9228 3556 11384 3564
rect 6536 3188 11384 3556
rect 6536 3172 7410 3188
rect 9228 3172 11384 3188
rect 14466 3576 15296 3946
rect 17228 3576 18058 3936
rect 14466 3558 18452 3576
rect 18778 3558 19324 8430
rect 14466 3144 19324 3558
rect 14486 3134 19324 3144
rect 19392 2012 19592 2212
rect -338 558 -138 758
rect -342 -3892 -142 -3692
<< via1 >>
rect 6076 5984 6770 6080
rect 8780 5984 9474 6080
rect 13930 5954 14624 6050
rect 16626 5960 17320 6056
<< metal2 >>
rect 6076 6080 6770 6090
rect 8780 6086 9474 6090
rect 6070 5984 6076 6036
rect 6070 5974 6770 5984
rect 8762 6080 9488 6086
rect 8762 5984 8780 6080
rect 9474 5984 9488 6080
rect 6070 5438 6762 5974
rect 6070 5404 6770 5438
rect 8762 5404 9488 5984
rect 13930 6050 14624 6060
rect 16626 6056 17320 6066
rect 13930 5944 14624 5954
rect 16604 5960 16626 6022
rect 17320 5960 17330 6022
rect 13930 5416 14622 5944
rect 16604 5416 17330 5960
rect 6070 5124 9488 5404
rect 13922 5152 17330 5416
rect 6070 3160 6770 5124
rect 13930 3196 14622 5152
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM1
timestamp 1752660100
transform 0 1 7751 -1 0 6037
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM2
timestamp 1752660100
transform 0 1 15607 -1 0 6011
box -2225 -2837 2225 2837
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM3
timestamp 1752660100
transform 1 0 15850 0 1 -1314
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM4
timestamp 1752660100
transform 1 0 18074 0 1 -1834
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM5
timestamp 1752660100
transform 1 0 19578 0 1 -1954
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM6
timestamp 1752660100
transform 1 0 14068 0 1 -1414
box -296 -610 296 610
use sky130_fd_pr__pfet_01v8_lvt_CYPNY8  XM7
timestamp 1752660100
transform 1 0 13009 0 1 2141
box -419 -519 419 519
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM8
timestamp 1752660100
transform 1 0 16895 0 1 479
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM9
timestamp 1752660100
transform 1 0 14991 0 1 839
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_CYPNY8  XM10
timestamp 1752660100
transform 1 0 14771 0 1 2241
box -419 -519 419 519
use sky130_fd_pr__pfet_01v8_lvt_6VJTDW  XM11
timestamp 1752660100
transform 1 0 22998 0 1 6790
box -936 -2332 946 2342
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR1
timestamp 1752660100
transform 1 0 17699 0 1 11860
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1752660100
transform 1 0 12029 0 1 -1564
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR3
timestamp 1752660100
transform 1 0 22129 0 1 -624
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_DBPYMX  XR4
timestamp 1752660100
transform 1 0 13271 0 1 12709
box -201 -889 201 889
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR5
timestamp 1752660100
transform 1 0 18881 0 1 11580
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR6
timestamp 1752660100
transform 1 0 21073 0 1 -624
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR7
timestamp 1752660100
transform 1 0 16177 0 1 12000
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_MAXMKG  XR8
timestamp 1752660100
transform 1 0 14573 0 1 12322
box -201 -742 201 742
<< labels >>
flabel metal1 19392 2012 19592 2212 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 -342 -3892 -142 -3692 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 -342 9256 -142 9456 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -338 558 -138 758 0 FreeSans 256 0 0 0 IN-
port 3 nsew
flabel metal1 -358 5854 -158 6054 0 FreeSans 256 0 0 0 IN+
port 4 nsew
<< end >>
