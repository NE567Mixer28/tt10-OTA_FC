magic
tech sky130A
magscale 1 2
timestamp 1770389351
<< metal3 >>
rect -6492 9332 -120 9360
rect -6492 3308 -204 9332
rect -140 3308 -120 9332
rect -6492 3280 -120 3308
rect 120 9332 6492 9360
rect 120 3308 6408 9332
rect 6472 3308 6492 9332
rect 120 3280 6492 3308
rect -6492 3012 -120 3040
rect -6492 -3012 -204 3012
rect -140 -3012 -120 3012
rect -6492 -3040 -120 -3012
rect 120 3012 6492 3040
rect 120 -3012 6408 3012
rect 6472 -3012 6492 3012
rect 120 -3040 6492 -3012
rect -6492 -3308 -120 -3280
rect -6492 -9332 -204 -3308
rect -140 -9332 -120 -3308
rect -6492 -9360 -120 -9332
rect 120 -3308 6492 -3280
rect 120 -9332 6408 -3308
rect 6472 -9332 6492 -3308
rect 120 -9360 6492 -9332
<< via3 >>
rect -204 3308 -140 9332
rect 6408 3308 6472 9332
rect -204 -3012 -140 3012
rect 6408 -3012 6472 3012
rect -204 -9332 -140 -3308
rect 6408 -9332 6472 -3308
<< mimcap >>
rect -6452 9280 -452 9320
rect -6452 3360 -6412 9280
rect -492 3360 -452 9280
rect -6452 3320 -452 3360
rect 160 9280 6160 9320
rect 160 3360 200 9280
rect 6120 3360 6160 9280
rect 160 3320 6160 3360
rect -6452 2960 -452 3000
rect -6452 -2960 -6412 2960
rect -492 -2960 -452 2960
rect -6452 -3000 -452 -2960
rect 160 2960 6160 3000
rect 160 -2960 200 2960
rect 6120 -2960 6160 2960
rect 160 -3000 6160 -2960
rect -6452 -3360 -452 -3320
rect -6452 -9280 -6412 -3360
rect -492 -9280 -452 -3360
rect -6452 -9320 -452 -9280
rect 160 -3360 6160 -3320
rect 160 -9280 200 -3360
rect 6120 -9280 6160 -3360
rect 160 -9320 6160 -9280
<< mimcapcontact >>
rect -6412 3360 -492 9280
rect 200 3360 6120 9280
rect -6412 -2960 -492 2960
rect 200 -2960 6120 2960
rect -6412 -9280 -492 -3360
rect 200 -9280 6120 -3360
<< metal4 >>
rect -3504 9281 -3400 9480
rect -224 9332 -120 9480
rect -6413 9280 -491 9281
rect -6413 3360 -6412 9280
rect -492 3360 -491 9280
rect -6413 3359 -491 3360
rect -3504 2961 -3400 3359
rect -224 3308 -204 9332
rect -140 3308 -120 9332
rect 3108 9281 3212 9480
rect 6388 9332 6492 9480
rect 199 9280 6121 9281
rect 199 3360 200 9280
rect 6120 3360 6121 9280
rect 199 3359 6121 3360
rect -224 3012 -120 3308
rect -6413 2960 -491 2961
rect -6413 -2960 -6412 2960
rect -492 -2960 -491 2960
rect -6413 -2961 -491 -2960
rect -3504 -3359 -3400 -2961
rect -224 -3012 -204 3012
rect -140 -3012 -120 3012
rect 3108 2961 3212 3359
rect 6388 3308 6408 9332
rect 6472 3308 6492 9332
rect 6388 3012 6492 3308
rect 199 2960 6121 2961
rect 199 -2960 200 2960
rect 6120 -2960 6121 2960
rect 199 -2961 6121 -2960
rect -224 -3308 -120 -3012
rect -6413 -3360 -491 -3359
rect -6413 -9280 -6412 -3360
rect -492 -9280 -491 -3360
rect -6413 -9281 -491 -9280
rect -3504 -9480 -3400 -9281
rect -224 -9332 -204 -3308
rect -140 -9332 -120 -3308
rect 3108 -3359 3212 -2961
rect 6388 -3012 6408 3012
rect 6472 -3012 6492 3012
rect 6388 -3308 6492 -3012
rect 199 -3360 6121 -3359
rect 199 -9280 200 -3360
rect 6120 -9280 6121 -3360
rect 199 -9281 6121 -9280
rect -224 -9480 -120 -9332
rect 3108 -9480 3212 -9281
rect 6388 -9332 6408 -3308
rect 6472 -9332 6492 -3308
rect 6388 -9480 6492 -9332
<< properties >>
string FIXED_BBOX 120 3280 6200 9360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
