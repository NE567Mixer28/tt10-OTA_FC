magic
tech sky130A
magscale 1 2
timestamp 1770543261
<< viali >>
rect 59806 3962 60014 4018
rect 4362 -990 4810 -906
rect 8348 -974 8798 -906
rect 12304 -1002 12744 -924
rect 75860 -936 76418 -872
rect 4368 -1316 4816 -1232
rect 65378 -1794 65886 -1738
rect 69154 -1760 69712 -1696
rect 73132 -1788 73690 -1724
rect -2320 -4962 -2234 -4742
rect -2334 -6710 -2248 -6490
rect 58388 -10762 58448 -10640
rect 64564 -10758 64608 -10630
rect 68398 -10766 68446 -10620
rect 74044 -10758 74146 -10622
rect 48224 -11160 48288 -10944
rect 60058 -11876 60094 -11754
rect 64180 -11922 64244 -11796
rect 70034 -11940 70090 -11808
rect 73440 -11948 73496 -11816
rect 51766 -13874 51850 -13710
rect 51748 -14930 51832 -14766
rect 51756 -16002 51840 -15838
rect 51770 -17190 51854 -17026
rect 4116 -22706 4522 -22660
rect 8296 -22706 8646 -22644
rect 12778 -22738 13126 -22670
rect 58288 -34148 58364 -33994
rect 58284 -35682 58360 -35528
rect 58318 -37092 58394 -36938
rect 58288 -38590 58364 -38436
rect 20154 -39604 20506 -39512
<< metal1 >>
rect -1576 15936 902 15940
rect -7928 15904 902 15936
rect -7928 15140 -1594 15904
rect -1604 15092 -1594 15140
rect -782 15136 902 15904
rect -782 15092 -772 15136
rect 15604 15128 31505 15902
rect -1586 15086 -782 15092
rect 46628 15058 63915 15832
rect 78291 15100 83645 15874
rect -1702 13486 402 13496
rect -1702 13230 -1688 13486
rect -1432 13230 402 13486
rect -1702 13196 402 13230
rect 15882 13468 18356 13496
rect 15882 13016 17812 13468
rect 17802 12982 17812 13016
rect 18346 12982 18356 13468
rect 29470 13398 31392 13430
rect 48862 13426 48872 13550
rect 29470 13142 29502 13398
rect 29758 13142 31392 13398
rect 29470 13112 31392 13142
rect 46906 12962 48872 13426
rect 49458 12962 49468 13550
rect 61674 13422 63604 13462
rect 61674 13166 61704 13422
rect 61960 13166 63604 13422
rect 61674 13122 63604 13166
rect 79058 13386 80716 13468
rect 79058 13000 80308 13386
rect 80694 13000 80716 13386
rect 79058 12988 80716 13000
rect 46906 12946 49414 12962
rect -266 9820 126 9822
rect -7906 9300 254 9820
rect 15889 9689 31898 9750
rect 15889 9271 16708 9689
rect 17126 9271 31898 9689
rect 15889 9228 31898 9271
rect 62611 9740 63861 9792
rect 62611 9364 62658 9740
rect 63034 9364 63861 9740
rect 62611 9270 63861 9364
rect 15889 8785 16411 9228
rect 47520 9094 47530 9146
rect 46994 8712 47530 9094
rect 47520 8526 47530 8712
rect 48150 9094 48160 9146
rect 48150 8712 53701 9094
rect 48150 8526 48160 8712
rect -2524 6645 -1875 6649
rect -952 6645 344 6722
rect -2524 6466 344 6645
rect -2524 -4323 -2345 6466
rect -952 6454 344 6466
rect -952 6278 -704 6454
rect -952 6238 -703 6278
rect -941 -981 -703 6238
rect 27398 6208 31826 6812
rect 15960 5634 19002 5966
rect 18670 4872 19002 5634
rect 16001 2696 16351 4687
rect 18486 4252 18496 4872
rect 19196 4252 19206 4872
rect 27398 4848 28002 6208
rect 46916 5564 48678 5896
rect 48346 5234 48678 5564
rect 27388 4244 27398 4848
rect 28002 4244 28012 4848
rect 48176 4716 48186 5234
rect 48736 4716 48746 5234
rect 16001 2346 30594 2696
rect 31064 2346 31074 2696
rect 33920 2368 33930 2874
rect 34260 2368 34270 2874
rect 46978 2826 47402 4654
rect 53319 4329 53701 8712
rect 79146 8754 83594 9136
rect 79146 8352 79528 8754
rect 79146 8011 79172 8352
rect 79162 7888 79172 8011
rect 79636 7888 79646 8352
rect 62585 6387 63507 6761
rect 53319 3947 59563 4329
rect 62585 4312 62959 6387
rect 79191 5533 81546 5959
rect 60270 4184 62959 4312
rect 60162 4068 60172 4184
rect 60480 4068 62959 4184
rect 59794 4018 60026 4024
rect 59794 3996 59806 4018
rect 59792 3962 59806 3996
rect 60014 3962 60026 4018
rect 59792 3956 60026 3962
rect 59792 3555 60006 3956
rect 60270 3938 62959 4068
rect 79184 3902 79512 4738
rect 59131 3341 59141 3555
rect 59355 3341 60006 3555
rect 79158 3546 79168 3902
rect 79524 3546 79534 3902
rect 46978 2402 62862 2826
rect 63306 2402 63316 2826
rect 66050 2472 66060 2934
rect 66350 2472 66360 2934
rect 46362 1116 46372 1786
rect 47102 1766 52296 1786
rect 47102 1154 51676 1766
rect 52296 1154 52306 1766
rect 58889 1514 59651 1541
rect 58889 1276 59128 1514
rect 59442 1276 59651 1514
rect 47102 1124 52296 1154
rect 47102 1116 47112 1124
rect 4358 -900 4814 178
rect 8350 -900 8802 128
rect 4350 -906 4822 -900
rect -941 -1010 1493 -981
rect 4350 -990 4362 -906
rect 4810 -990 4822 -906
rect 8336 -906 8810 -900
rect 8336 -974 8348 -906
rect 8798 -974 8810 -906
rect 12308 -918 12750 82
rect 15153 4 31629 766
rect 58889 696 59651 1276
rect 46628 -66 63671 696
rect 27406 -832 27416 -816
rect 8336 -980 8810 -974
rect 12292 -924 12756 -918
rect 8350 -982 8802 -980
rect 4350 -996 4822 -990
rect -941 -1216 3290 -1010
rect 5758 -1182 7214 -1008
rect 9810 -1190 11334 -996
rect 12292 -1002 12304 -924
rect 12744 -1002 12756 -924
rect 12292 -1008 12756 -1002
rect 16698 -1016 16708 -924
rect 13838 -1182 16708 -1016
rect -941 -1219 1493 -1216
rect 4356 -1232 4828 -1226
rect 4356 -1316 4368 -1232
rect 4816 -1316 4828 -1232
rect 4356 -1322 4828 -1316
rect -2518 -4560 -2352 -4323
rect -2326 -4738 -2228 -4730
rect 4474 -4738 4694 -1322
rect 16698 -1350 16708 -1182
rect 17132 -1350 17142 -924
rect 18585 -1485 18595 -1111
rect 18969 -1485 18979 -1111
rect 27396 -1420 27416 -832
rect 28020 -832 28030 -816
rect 28020 -1420 46414 -832
rect 27396 -1440 46414 -1420
rect 47022 -1440 47032 -832
rect 18595 -4067 18969 -1485
rect 48253 -1521 48263 -1147
rect 48637 -1521 48647 -1147
rect 48263 -4067 48637 -1521
rect 65374 -1732 65890 78
rect 69174 -1690 69690 102
rect 69142 -1696 69724 -1690
rect 63096 -2062 63106 -1734
rect 63434 -1744 63444 -1734
rect 65366 -1738 65898 -1732
rect 63434 -2062 64338 -1744
rect 65366 -1794 65378 -1738
rect 65886 -1794 65898 -1738
rect 65366 -1800 65898 -1794
rect 63108 -2072 64338 -2062
rect 66784 -2170 68252 -1730
rect 69142 -1760 69154 -1696
rect 69712 -1760 69724 -1696
rect 69142 -1766 69724 -1760
rect 69174 -1770 69690 -1766
rect 70748 -2078 72082 -1678
rect 73114 -1718 73688 126
rect 75868 -866 76426 156
rect 75848 -872 76430 -866
rect 75848 -936 75860 -872
rect 76418 -936 76430 -872
rect 75848 -942 76430 -936
rect 73114 -1724 73702 -1718
rect 73114 -1782 73132 -1724
rect 73120 -1788 73132 -1782
rect 73690 -1788 73702 -1724
rect 73120 -1794 73702 -1788
rect 74550 -1970 74884 -996
rect 77190 -1620 77532 -938
rect 77112 -2058 77122 -1620
rect 77668 -2058 77678 -1620
rect 18550 -4441 59307 -4067
rect -2326 -4742 4694 -4738
rect -2326 -4962 -2320 -4742
rect -2234 -4958 4694 -4742
rect -2234 -4962 -2228 -4958
rect -2326 -4974 -2228 -4962
rect -3788 -5620 -3411 -5618
rect -2518 -5620 -2356 -5064
rect -3788 -5776 -2356 -5620
rect -3790 -5804 -2356 -5776
rect -3790 -5884 -3410 -5804
rect -3790 -6058 -3404 -5884
rect -3790 -6680 -3410 -6058
rect -2518 -6372 -2356 -5804
rect -2340 -6490 -2242 -6478
rect -7886 -12884 -7026 -12368
rect -7036 -12898 -7026 -12884
rect -6338 -12898 -6328 -12368
rect -3782 -33342 -3415 -6680
rect -2340 -6710 -2334 -6490
rect -2248 -6494 -2242 -6490
rect -1912 -6494 -1692 -4958
rect -2248 -6710 -1692 -6494
rect -2340 -6722 -2242 -6710
rect -1912 -6712 -1692 -6710
rect -2554 -15577 -2375 -6786
rect -1288 -7050 -1278 -6246
rect -474 -7050 938 -6246
rect 15337 -7058 31489 -6284
rect 46459 -7132 56701 -6358
rect 46871 -7770 46881 -7739
rect 62 -7970 476 -7913
rect 48 -8226 58 -7970
rect 314 -8226 476 -7970
rect 62 -9002 476 -8226
rect 46804 -8173 46881 -7770
rect 47315 -8173 47325 -7739
rect 15702 -8719 17895 -8690
rect 15702 -9153 17435 -8719
rect 17869 -9153 17895 -8719
rect 30163 -8756 31362 -8662
rect 30163 -9012 30270 -8756
rect 30526 -9012 31362 -8756
rect 30163 -9076 31362 -9012
rect 15702 -9176 17895 -9153
rect 46804 -9244 47284 -8173
rect 48906 -8228 48916 -7896
rect 49248 -8228 49258 -7896
rect 48916 -9249 49248 -8228
rect 55927 -8633 56701 -7132
rect 58933 -7220 59307 -4441
rect 58933 -7256 68264 -7220
rect 58933 -7594 67944 -7256
rect 67934 -7648 67944 -7594
rect 68300 -7648 68310 -7256
rect 47944 -9296 48276 -9276
rect 48805 -9296 52320 -9249
rect 47944 -9628 52320 -9296
rect 55927 -9407 72535 -8633
rect 73566 -9108 73576 -8732
rect 73952 -9108 73962 -8732
rect 47944 -10714 48276 -9628
rect 48805 -9651 52320 -9628
rect 48218 -10936 48294 -10932
rect 48218 -10944 49698 -10936
rect 48218 -11160 48224 -10944
rect 48288 -11160 49698 -10944
rect 48218 -11172 49698 -11160
rect 45764 -11629 48167 -11263
rect 48224 -11298 49698 -11172
rect -731 -12888 -721 -12366
rect -199 -12888 582 -12366
rect 29803 -12931 31067 -12549
rect 19335 -13022 19345 -13021
rect 15725 -13404 19345 -13022
rect 19335 -13407 19345 -13404
rect 19731 -13022 19741 -13021
rect 29803 -13022 30185 -12931
rect 19731 -13404 30185 -13022
rect 47597 -13096 47607 -12965
rect 19731 -13407 19741 -13404
rect 46892 -13478 47607 -13096
rect 47597 -13627 47607 -13478
rect 48269 -13627 48279 -12965
rect 49336 -13917 49698 -11298
rect 51760 -13710 51856 -13698
rect 51074 -13714 51512 -13710
rect 51760 -13714 51766 -13710
rect 51074 -13870 51766 -13714
rect 51074 -13917 51512 -13870
rect 51760 -13874 51766 -13870
rect 51850 -13874 51856 -13710
rect 51918 -13820 52320 -9651
rect 56520 -10712 56790 -9407
rect 57958 -9756 58226 -9744
rect 57958 -9996 57974 -9756
rect 58232 -9996 58242 -9756
rect 57958 -10653 58226 -9996
rect 58382 -10638 58454 -10628
rect 58382 -10640 59846 -10638
rect 57939 -11095 58237 -10653
rect 58382 -10762 58388 -10640
rect 58448 -10762 59846 -10640
rect 62714 -10704 62984 -9407
rect 64098 -10210 64108 -9868
rect 64444 -10210 64454 -9868
rect 64108 -10704 64430 -10210
rect 64558 -10630 64614 -10618
rect 58382 -10770 59846 -10762
rect 58382 -10774 58454 -10770
rect 56580 -11393 58237 -11095
rect 56580 -11848 56878 -11393
rect 59714 -11750 59846 -10770
rect 64123 -11105 64421 -10704
rect 64558 -10758 64564 -10630
rect 64608 -10634 64614 -10630
rect 64608 -10744 65156 -10634
rect 66560 -10704 66830 -9407
rect 67932 -10188 67942 -9886
rect 68270 -10188 68280 -9886
rect 67950 -10671 68248 -10188
rect 68410 -10608 69882 -10604
rect 67947 -10726 68248 -10671
rect 68392 -10620 69882 -10608
rect 64608 -10758 64614 -10744
rect 64558 -10770 64614 -10758
rect 62734 -11403 64421 -11105
rect 60052 -11750 60100 -11742
rect 59642 -11754 60210 -11750
rect 59642 -11876 60058 -11754
rect 60094 -11876 60210 -11754
rect 62734 -11784 63032 -11403
rect 59642 -13147 60210 -11876
rect 62732 -11858 63032 -11784
rect 64174 -11792 64250 -11784
rect 63780 -11796 64328 -11792
rect 62732 -12414 63030 -11858
rect 63780 -11922 64180 -11796
rect 64244 -11922 64328 -11796
rect 62662 -12712 62672 -12414
rect 63158 -12712 63168 -12414
rect 63780 -13147 64328 -11922
rect 65042 -13147 65146 -10744
rect 66546 -11149 66844 -11139
rect 67947 -11149 68245 -10726
rect 68392 -10766 68398 -10620
rect 68446 -10766 69882 -10620
rect 72206 -10690 72476 -9407
rect 73596 -10683 73886 -9108
rect 74241 -10604 74432 -10602
rect 74038 -10612 74152 -10610
rect 74202 -10612 74432 -10604
rect 74038 -10622 74432 -10612
rect 68392 -10778 69882 -10766
rect 73596 -10770 73895 -10683
rect 74038 -10758 74044 -10622
rect 74146 -10758 74432 -10622
rect 74038 -10770 74432 -10758
rect 68410 -10784 69882 -10778
rect 66546 -11447 68245 -11149
rect 66546 -11892 66844 -11447
rect 69704 -11798 69881 -10784
rect 73597 -11135 73895 -10770
rect 74082 -10772 74432 -10770
rect 74202 -10808 74432 -10772
rect 72276 -11433 73895 -11135
rect 70028 -11798 70096 -11796
rect 69608 -11808 70116 -11798
rect 66546 -12386 66842 -11892
rect 69608 -11940 70034 -11808
rect 70090 -11940 70116 -11808
rect 72276 -11892 72574 -11433
rect 73434 -11816 73502 -11804
rect 73434 -11818 73440 -11816
rect 66536 -12598 66546 -12386
rect 66848 -12598 66858 -12386
rect 69608 -13147 70116 -11940
rect 72282 -12370 72572 -11892
rect 73024 -11948 73440 -11818
rect 73496 -11948 73502 -11816
rect 73024 -11960 73502 -11948
rect 72168 -12820 72178 -12370
rect 72618 -12820 72628 -12370
rect 73024 -13147 73470 -11960
rect 74241 -13147 74432 -10808
rect 78655 -13147 79417 781
rect 81120 -7287 81546 5533
rect 81120 -7601 81181 -7287
rect 81495 -7601 81546 -7287
rect 81120 -7682 81546 -7601
rect 51760 -13886 51856 -13874
rect 49336 -14279 51512 -13917
rect 54624 -14147 54942 -13722
rect 51074 -14770 51512 -14279
rect 51939 -14465 54942 -14147
rect 59373 -13909 79417 -13147
rect 51742 -14766 51838 -14754
rect 51742 -14770 51748 -14766
rect 51074 -14926 51748 -14770
rect -960 -15472 18 -15432
rect -960 -15577 292 -15472
rect -2554 -15756 292 -15577
rect -962 -15757 292 -15756
rect -960 -15832 292 -15757
rect -960 -22568 -722 -15832
rect -694 -15834 292 -15832
rect 28682 -15982 31724 -15378
rect 51074 -15828 51512 -14926
rect 51742 -14930 51748 -14926
rect 51832 -14930 51838 -14766
rect 51939 -14895 52257 -14465
rect 51742 -14942 51838 -14930
rect 54610 -15138 54888 -14832
rect 51987 -15416 54888 -15138
rect 51750 -15828 51846 -15826
rect 51074 -15838 51846 -15828
rect 16002 -16312 17722 -16220
rect 16002 -16552 17428 -16312
rect 17418 -16640 17428 -16552
rect 17756 -16640 17766 -16312
rect 16036 -18229 16448 -17482
rect 16025 -18643 16035 -18229
rect 16449 -18643 16459 -18229
rect 28682 -18338 29286 -15982
rect 51074 -15984 51756 -15838
rect 46888 -16340 48768 -16294
rect 46888 -16626 48444 -16340
rect 48434 -16668 48444 -16626
rect 48772 -16668 48782 -16340
rect 51074 -17016 51512 -15984
rect 51750 -16002 51756 -15984
rect 51840 -16002 51846 -15838
rect 51987 -15957 52265 -15416
rect 51750 -16014 51846 -16002
rect 54582 -16366 54874 -15818
rect 51980 -16658 54874 -16366
rect 51764 -17016 51860 -17014
rect 51074 -17026 51860 -17016
rect 51074 -17172 51770 -17026
rect 16036 -18650 16448 -18643
rect 28672 -18942 28682 -18338
rect 29286 -18942 29296 -18338
rect 46888 -18397 47264 -17522
rect 46888 -18739 46905 -18397
rect 47247 -18739 47264 -18397
rect 51074 -18057 51512 -17172
rect 51764 -17190 51770 -17172
rect 51854 -17190 51860 -17026
rect 51980 -17156 52272 -16658
rect 51764 -17202 51860 -17190
rect 54624 -17288 56802 -16942
rect 56456 -17543 56802 -17288
rect 56456 -17889 57449 -17543
rect 57795 -17889 57805 -17543
rect 51074 -18495 53013 -18057
rect 46888 -18798 47264 -18739
rect 33852 -19690 33862 -19200
rect 34170 -19690 34180 -19200
rect -962 -22706 -716 -22568
rect 4124 -22654 4514 -22092
rect 8302 -22638 8654 -22070
rect 8284 -22644 8658 -22638
rect 4104 -22660 4534 -22654
rect 4104 -22706 4116 -22660
rect 4522 -22706 4534 -22660
rect -976 -22932 2948 -22706
rect 4104 -22712 4534 -22706
rect 8284 -22706 8296 -22644
rect 8646 -22706 8658 -22644
rect 12774 -22664 13134 -22008
rect 15411 -22182 31889 -21420
rect 52575 -21494 53013 -18495
rect 59373 -21494 60135 -13909
rect 68047 -15515 71945 -15009
rect 72451 -15515 72461 -15009
rect 68047 -16101 68553 -15515
rect 46309 -22256 60135 -21494
rect 61341 -16607 68553 -16101
rect 8284 -22712 8658 -22706
rect 12766 -22670 13138 -22664
rect 5546 -22922 7314 -22720
rect 12766 -22738 12778 -22670
rect 13126 -22738 13138 -22670
rect 9754 -22940 11832 -22738
rect 12766 -22744 13138 -22738
rect 14052 -23438 14440 -22800
rect 14052 -23826 16802 -23438
rect 17190 -23826 17200 -23438
rect 23162 -25358 23172 -24766
rect 23764 -24818 23774 -24766
rect 57624 -24818 57634 -24746
rect 23764 -25358 57634 -24818
rect 57624 -25510 57634 -25358
rect 58480 -25510 58490 -24746
rect 21816 -26678 21826 -26098
rect 22594 -26112 22604 -26098
rect 24846 -26112 24856 -26098
rect 22594 -26678 24856 -26112
rect 21826 -26704 24856 -26678
rect 25798 -26704 25808 -26098
rect -1992 -27294 1066 -27222
rect -1992 -28026 -1856 -27294
rect -1866 -28101 -1856 -28026
rect -1049 -28026 1066 -27294
rect -1049 -28101 -1039 -28026
rect 15169 -28034 31487 -27260
rect -88 -28932 326 -28903
rect -130 -29188 -120 -28932
rect 136 -29188 326 -28932
rect 14174 -29078 14184 -28602
rect 14978 -29078 14988 -28602
rect -88 -29978 326 -29188
rect 23225 -29617 23235 -29095
rect 23757 -29617 23767 -29095
rect 15768 -30146 16872 -29666
rect 17352 -30146 17362 -29666
rect -3782 -33657 204 -33342
rect -3774 -33864 204 -33657
rect 23235 -33346 23757 -29617
rect 29451 -29654 31288 -29568
rect 29451 -29910 29476 -29654
rect 29732 -29910 31288 -29654
rect 48224 -29670 48234 -29576
rect 29451 -29982 31288 -29910
rect 46514 -30060 48234 -29670
rect 48718 -29610 48728 -29576
rect 61341 -29610 61847 -16607
rect 48718 -30060 61847 -29610
rect 46514 -30116 61847 -30060
rect 46514 -30156 48719 -30116
rect 55084 -32322 55094 -31772
rect 55696 -32322 55706 -31772
rect 23235 -33868 31394 -33346
rect 16588 -33987 16598 -33876
rect 16573 -33998 16598 -33987
rect 15856 -34380 16598 -33998
rect 16573 -34396 16598 -34380
rect 17118 -33987 17128 -33876
rect 17118 -34396 17187 -33987
rect 46805 -34384 53067 -34002
rect 55188 -34142 55522 -32322
rect 58282 -33994 58370 -33982
rect 58616 -33994 59128 -33990
rect 16573 -35449 17187 -34396
rect 16573 -36063 19264 -35449
rect -7060 -36884 -7050 -36280
rect -6446 -36884 688 -36280
rect 15964 -37510 17298 -37262
rect 15850 -39086 16184 -38426
rect 15850 -39313 15938 -39086
rect 15928 -39326 15938 -39313
rect 16178 -39326 16188 -39086
rect 17050 -40426 17298 -37510
rect 18650 -38594 19264 -36063
rect 28232 -36816 28242 -36128
rect 28982 -36288 28992 -36128
rect 28982 -36816 31468 -36288
rect 28276 -36884 31468 -36816
rect 18650 -39208 19776 -38594
rect 28276 -38602 28872 -36884
rect 47882 -37200 47892 -37184
rect 20800 -39198 28872 -38602
rect 29988 -37364 30236 -37332
rect 33906 -37364 34090 -37348
rect 29988 -37548 34090 -37364
rect 46804 -37512 47892 -37200
rect 48220 -37512 48230 -37184
rect 46804 -37532 48214 -37512
rect 20146 -39506 20522 -39500
rect 20142 -39512 20522 -39506
rect 20142 -39604 20154 -39512
rect 20506 -39604 20522 -39512
rect 20142 -39610 20522 -39604
rect 18534 -40426 18544 -40340
rect 17050 -40674 18544 -40426
rect 18534 -40818 18544 -40674
rect 19060 -40818 19070 -40340
rect -8058 -43160 901 -42394
rect 20146 -42396 20522 -39610
rect 21656 -40818 21666 -40346
rect 22212 -40426 22222 -40346
rect 29988 -40426 30236 -37548
rect 33906 -38204 34090 -37548
rect 52685 -38146 53067 -34384
rect 55210 -37024 55572 -35598
rect 57810 -35636 58134 -34046
rect 58282 -34148 58288 -33994
rect 58364 -34148 59128 -33994
rect 58282 -34160 58370 -34148
rect 58278 -35524 58366 -35516
rect 58616 -35524 59128 -34148
rect 58278 -35528 59128 -35524
rect 58278 -35682 58284 -35528
rect 58360 -35678 59128 -35528
rect 58360 -35682 58366 -35678
rect 58278 -35694 58366 -35682
rect 58616 -36922 59128 -35678
rect 58326 -36926 59128 -36922
rect 58312 -36938 59128 -36926
rect 46812 -38461 49929 -38430
rect 46812 -38764 49589 -38461
rect 49579 -38803 49589 -38764
rect 49931 -38803 49941 -38461
rect 52516 -38854 52526 -38146
rect 53192 -38375 53202 -38146
rect 53192 -38757 55371 -38375
rect 57862 -38554 58134 -36986
rect 58312 -37092 58318 -36938
rect 58394 -37076 59128 -36938
rect 58394 -37092 58400 -37076
rect 58312 -37104 58400 -37092
rect 58282 -38436 58370 -38424
rect 58616 -38436 59128 -37076
rect 58282 -38590 58288 -38436
rect 58364 -38590 59128 -38436
rect 58282 -38602 58370 -38590
rect 53192 -38854 53202 -38757
rect 22212 -40674 30236 -40426
rect 33786 -40668 33796 -40202
rect 34104 -40668 34114 -40202
rect 22212 -40818 22222 -40674
rect 15411 -43158 31457 -42396
rect 58616 -42400 59128 -38590
rect 78655 -42400 79417 -13909
rect 80444 -17382 83594 -17368
rect 80404 -18100 80414 -17382
rect 81016 -18100 83594 -17382
rect 80854 -19874 83578 -19860
rect 80316 -20592 80326 -19874
rect 80928 -20592 83578 -19874
rect 80404 -25456 80414 -24738
rect 81016 -25456 83550 -24738
rect 80516 -25544 83550 -25456
rect 46099 -43162 79417 -42400
<< via1 >>
rect -1594 15092 -782 15904
rect -1688 13230 -1432 13486
rect 17812 12982 18346 13468
rect 29502 13142 29758 13398
rect 48872 12962 49458 13550
rect 61704 13166 61960 13422
rect 80308 13000 80694 13386
rect 16708 9271 17126 9689
rect 62658 9364 63034 9740
rect 47530 8526 48150 9146
rect 18496 4252 19196 4872
rect 27398 4244 28002 4848
rect 48186 4716 48736 5234
rect 30594 2346 31064 2696
rect 33930 2368 34260 2874
rect 79172 7888 79636 8352
rect 60172 4068 60480 4184
rect 59141 3341 59355 3555
rect 79168 3546 79524 3902
rect 62862 2402 63306 2826
rect 66060 2472 66350 2934
rect 46372 1116 47102 1786
rect 51676 1154 52296 1766
rect 59128 1276 59442 1514
rect 16708 -1350 17132 -924
rect 18595 -1485 18969 -1111
rect 27416 -1420 28020 -816
rect 46414 -1440 47022 -832
rect 48263 -1521 48637 -1147
rect 63106 -2062 63434 -1734
rect 77122 -2058 77668 -1620
rect -7026 -12898 -6338 -12368
rect -1278 -7050 -474 -6246
rect 58 -8226 314 -7970
rect 46881 -8173 47315 -7739
rect 17435 -9153 17869 -8719
rect 30270 -9012 30526 -8756
rect 48916 -8228 49248 -7896
rect 67944 -7648 68300 -7256
rect 73576 -9108 73952 -8732
rect -721 -12888 -199 -12366
rect 19345 -13407 19731 -13021
rect 47607 -13627 48269 -12965
rect 57974 -9996 58232 -9756
rect 64108 -10210 64444 -9868
rect 67942 -10188 68270 -9886
rect 62672 -12712 63158 -12414
rect 66546 -12598 66848 -12386
rect 72178 -12820 72618 -12370
rect 81181 -7601 81495 -7287
rect 17428 -16640 17756 -16312
rect 16035 -18643 16449 -18229
rect 48444 -16668 48772 -16340
rect 28682 -18942 29286 -18338
rect 46905 -18739 47247 -18397
rect 57449 -17889 57795 -17543
rect 33862 -19690 34170 -19200
rect 71945 -15515 72451 -15009
rect 16802 -23826 17190 -23438
rect 23172 -25358 23764 -24766
rect 57634 -25510 58480 -24746
rect 21826 -26678 22594 -26098
rect 24856 -26704 25798 -26098
rect -1856 -28101 -1049 -27294
rect -120 -29188 136 -28932
rect 14184 -29078 14978 -28602
rect 23235 -29617 23757 -29095
rect 16872 -30146 17352 -29666
rect 29476 -29910 29732 -29654
rect 48234 -30060 48718 -29576
rect 55094 -32322 55696 -31772
rect 16598 -34396 17118 -33876
rect -7050 -36884 -6446 -36280
rect 15938 -39326 16178 -39086
rect 28242 -36816 28982 -36128
rect 47892 -37512 48220 -37184
rect 18544 -40818 19060 -40340
rect 21666 -40818 22212 -40346
rect 49589 -38803 49931 -38461
rect 52526 -38854 53192 -38146
rect 33796 -40668 34104 -40202
rect 80414 -18100 81016 -17382
rect 80326 -20592 80928 -19874
rect 80414 -25456 81016 -24738
<< metal2 >>
rect -1594 15904 -782 15914
rect -4198 15092 -1594 15904
rect -782 15092 -776 15904
rect -4198 -1666 -3386 15092
rect -1594 15082 -782 15092
rect 48872 13550 49458 13560
rect -1688 13486 -1432 13496
rect -1688 -446 -1432 13230
rect 17812 13468 18346 13478
rect 17812 12972 18346 12982
rect 29502 13398 29758 13408
rect 16708 9689 17126 9699
rect -1688 -702 1068 -446
rect -5658 -2478 -463 -1666
rect -7026 -12368 -6338 -12358
rect -7026 -12908 -6338 -12898
rect -5655 -27294 -4848 -2478
rect -1275 -5899 -463 -2478
rect 812 -5188 1068 -702
rect 16708 -914 17126 9271
rect 18496 4872 19196 4882
rect 18496 4242 19196 4252
rect 27398 4848 28002 4858
rect 16708 -924 17132 -914
rect 16708 -1360 17132 -1350
rect 18584 -1111 18998 4242
rect 27398 4234 28002 4244
rect 18584 -1460 18595 -1111
rect 18969 -1460 18998 -1111
rect 27416 -806 27964 4234
rect 27416 -816 28020 -806
rect 27416 -1430 28020 -1420
rect 18595 -1495 18969 -1485
rect 29502 -5188 29758 13142
rect 48872 12952 49458 12962
rect 61704 13422 61960 13432
rect 47530 9146 48150 9156
rect 47530 7690 48150 8526
rect 47530 7070 52266 7690
rect 48186 5234 48736 5244
rect 48186 4706 48736 4716
rect 33930 2874 34260 2884
rect 30594 2696 31064 2706
rect 31064 2398 33930 2642
rect 33930 2358 34260 2368
rect 30594 2336 31064 2346
rect 46372 1786 47102 1796
rect 46372 1106 47102 1116
rect 46412 -832 47042 1106
rect 46412 -1440 46414 -832
rect 47022 -1440 47042 -832
rect 48260 -1147 48650 4706
rect 51646 1776 52266 7070
rect 60178 4194 60508 4210
rect 60172 4184 60508 4194
rect 60480 4068 60508 4184
rect 60172 4058 60508 4068
rect 59141 3555 59355 3565
rect 59134 3341 59141 3534
rect 59355 3341 59408 3534
rect 51646 1766 52296 1776
rect 51646 1196 51676 1766
rect 59134 1524 59408 3341
rect 60178 1714 60508 4058
rect 60178 1704 60534 1714
rect 59128 1514 59442 1524
rect 60178 1454 60186 1704
rect 60186 1372 60534 1382
rect 59128 1266 59442 1276
rect 51676 1144 52296 1154
rect 61704 -1076 61960 13166
rect 80308 13386 80694 13396
rect 80694 13000 80697 13361
rect 80308 12990 80697 13000
rect 62658 9740 63034 9750
rect 62658 9354 63034 9364
rect 79172 8352 79636 8362
rect 79172 7878 79636 7888
rect 80311 7485 80697 12990
rect 80311 7099 82585 7485
rect 79168 3902 79524 3912
rect 66060 2934 66350 2944
rect 62862 2826 63306 2836
rect 63306 2476 66060 2756
rect 66060 2462 66350 2472
rect 62862 2392 63306 2402
rect 79168 2290 79524 3546
rect 79168 1934 80458 2290
rect 46414 -1450 47022 -1440
rect 48260 -1506 48263 -1147
rect 48637 -1506 48650 -1147
rect 57964 -1332 61960 -1076
rect 48263 -1531 48637 -1521
rect 57964 -5188 58220 -1332
rect 77122 -1620 77668 -1610
rect 63106 -1734 63434 -1724
rect 63106 -2072 63434 -2062
rect 77122 -2068 77668 -2058
rect 614 -5444 58220 -5188
rect -1270 -6236 -468 -5899
rect -1278 -6246 -468 -6236
rect -474 -7028 -468 -6246
rect -1278 -7060 -474 -7050
rect 614 -7352 870 -5444
rect 58 -7490 870 -7352
rect -1526 -7608 870 -7490
rect -1526 -7746 314 -7608
rect -1526 -26258 -1270 -7746
rect 58 -7970 314 -7746
rect 58 -8236 314 -8226
rect 17435 -8719 17869 -8709
rect 29454 -8756 29710 -5444
rect 46881 -7739 47315 -7729
rect 46881 -8183 47315 -8173
rect 48916 -7896 49248 -7886
rect 48916 -8238 49248 -8228
rect 30270 -8756 30526 -8746
rect 29454 -9012 30270 -8756
rect 30270 -9022 30526 -9012
rect 17435 -9163 17869 -9153
rect 57964 -9746 58220 -5444
rect 80102 -5642 80458 1934
rect 64114 -5998 80458 -5642
rect 64114 -7302 64470 -5998
rect 67944 -7256 68300 -7246
rect 64094 -7446 64470 -7302
rect 57964 -9756 58232 -9746
rect 57964 -9996 57974 -9756
rect 57964 -10006 58232 -9996
rect 64094 -9868 64450 -7446
rect 57964 -10012 58220 -10006
rect 64094 -10210 64108 -9868
rect 64444 -10210 64450 -9868
rect 67942 -7648 67944 -7287
rect 81181 -7287 81495 -7277
rect 68300 -7601 81181 -7287
rect 81181 -7611 81495 -7601
rect 67942 -7658 68300 -7648
rect 67942 -9876 68256 -7658
rect 73546 -8634 74008 -8624
rect 82199 -8732 82585 7099
rect 74008 -9118 82585 -8732
rect 73546 -9162 74008 -9152
rect 67942 -9886 68270 -9876
rect 67942 -10198 68270 -10188
rect 64094 -10216 64450 -10210
rect 64108 -10220 64444 -10216
rect -721 -12366 -199 -12356
rect 72178 -12370 72618 -12360
rect 66546 -12386 66848 -12376
rect 62672 -12414 63158 -12404
rect 66546 -12608 66848 -12598
rect 62672 -12722 63158 -12712
rect -721 -12898 -199 -12888
rect 47607 -12965 48269 -12955
rect 19345 -13021 19731 -13011
rect 19345 -13417 19731 -13407
rect 47607 -13637 48269 -13627
rect 17428 -16312 17756 -16302
rect 17428 -16650 17756 -16640
rect 48444 -16340 48772 -16330
rect 48444 -16678 48772 -16668
rect 57449 -17543 57795 -17533
rect 57449 -17899 57795 -17889
rect 16035 -18229 16449 -18219
rect 16035 -20361 16449 -18643
rect 28682 -18338 29286 -18328
rect 28682 -18952 29286 -18942
rect 46905 -18397 47247 -18387
rect 33862 -19200 34170 -19190
rect 31153 -19690 33862 -19466
rect 31153 -19700 34170 -19690
rect 31153 -19880 34162 -19700
rect 31153 -20361 31567 -19880
rect 16035 -20775 31567 -20361
rect 46905 -20413 47247 -18739
rect 62714 -20413 63056 -12722
rect 71954 -12820 72178 -12576
rect 71954 -12830 72618 -12820
rect 71954 -14999 72480 -12830
rect 71945 -15009 72480 -14999
rect 72451 -15466 72480 -15009
rect 71945 -15525 72451 -15515
rect 80414 -17382 81016 -17372
rect 80414 -18110 81016 -18100
rect 46905 -20755 63056 -20413
rect 80326 -19874 80928 -19864
rect 80326 -20602 80928 -20592
rect 16802 -23438 17190 -23428
rect 16802 -23836 17190 -23826
rect 23172 -24766 23764 -24756
rect 21826 -26098 22594 -26088
rect -1526 -26514 21826 -26258
rect -1856 -27294 -1049 -27284
rect -5655 -28101 -1856 -27294
rect -1856 -28111 -1049 -28101
rect -120 -28932 136 -26514
rect 21826 -26688 22594 -26678
rect 14184 -28602 14978 -28592
rect 14978 -29078 19486 -28602
rect 14184 -29122 19486 -29078
rect 23172 -29095 23764 -25358
rect 24856 -26098 25798 -26088
rect 25798 -26514 29732 -26258
rect 24856 -26714 25798 -26704
rect -120 -29198 136 -29188
rect 16872 -29666 17352 -29656
rect 16872 -30156 17352 -30146
rect 16598 -33876 17118 -33866
rect 18908 -33876 19428 -29122
rect 23172 -29478 23235 -29095
rect 23757 -29478 23764 -29095
rect 23235 -29627 23757 -29617
rect 29476 -29654 29732 -26514
rect 29476 -29920 29732 -29910
rect 48234 -29576 48718 -29566
rect 48234 -30070 48718 -30060
rect 17118 -34396 19428 -33876
rect 16598 -34406 17118 -34396
rect 28242 -36128 28982 -36118
rect -7370 -36160 -6216 -36150
rect 28242 -36826 28982 -36816
rect -7370 -36950 -6216 -36940
rect 47892 -37184 48220 -37174
rect 47892 -37522 48220 -37512
rect 49589 -38461 49931 -20755
rect 57634 -24746 58480 -24736
rect 80414 -24738 81016 -24728
rect 58480 -25412 80414 -24776
rect 80414 -25466 81016 -25456
rect 57634 -25520 58480 -25510
rect 62453 -27949 63147 -27939
rect 58939 -28643 62453 -27949
rect 55094 -31772 55696 -31762
rect 55094 -32332 55696 -32322
rect 58939 -32385 59633 -28643
rect 62453 -28653 63147 -28643
rect 58939 -33079 62525 -32385
rect 49589 -38813 49931 -38803
rect 52526 -38146 53192 -38136
rect 53192 -38854 53220 -38188
rect 15938 -39086 16178 -39076
rect 15938 -41560 16178 -39326
rect 52526 -39692 53220 -38854
rect 61831 -39692 62525 -33079
rect 33796 -40202 34104 -40192
rect 18544 -40340 19060 -40330
rect 18398 -40700 18544 -40428
rect 21666 -40346 22212 -40336
rect 19060 -40700 21666 -40428
rect 18544 -40828 19060 -40818
rect 21666 -40828 22212 -40818
rect 30928 -40664 33796 -40424
rect 30928 -41560 31168 -40664
rect 52526 -40386 62525 -39692
rect 33796 -40678 34104 -40668
rect 15938 -41800 31168 -41560
<< via2 >>
rect 17812 12982 18346 13468
rect -7026 -12898 -6338 -12368
rect 48872 12962 49458 13550
rect 60186 1382 60534 1704
rect 62658 9364 63034 9740
rect 79172 7888 79636 8352
rect 63106 -2062 63434 -1734
rect 77122 -2058 77668 -1620
rect 17435 -9153 17869 -8719
rect 46881 -8173 47315 -7739
rect 48916 -8228 49248 -7896
rect 73546 -8732 74008 -8634
rect 73546 -9108 73576 -8732
rect 73576 -9108 73952 -8732
rect 73952 -9108 74008 -8732
rect 73546 -9152 74008 -9108
rect -721 -12888 -199 -12366
rect 66546 -12598 66848 -12386
rect 19345 -13407 19731 -13021
rect 47607 -13627 48269 -12965
rect 17428 -16640 17756 -16312
rect 48444 -16668 48772 -16340
rect 57449 -17889 57795 -17543
rect 28682 -18942 29286 -18338
rect 80414 -18100 81016 -17382
rect 80326 -20592 80928 -19874
rect 16802 -23826 17190 -23438
rect 14184 -29078 14978 -28602
rect 16872 -30146 17352 -29666
rect 48234 -30060 48718 -29576
rect -7370 -36280 -6216 -36160
rect -7370 -36884 -7050 -36280
rect -7050 -36884 -6446 -36280
rect -6446 -36884 -6216 -36280
rect 28242 -36816 28982 -36128
rect -7370 -36940 -6216 -36884
rect 47892 -37512 48220 -37184
rect 62453 -28643 63147 -27949
rect 55094 -32322 55696 -31772
<< metal3 >>
rect 48862 13550 49468 13555
rect 17837 13473 18271 13501
rect 17802 13468 18356 13473
rect 17802 12982 17812 13468
rect 18346 12982 18356 13468
rect 17802 12977 18356 12982
rect 17837 7605 18271 12977
rect 48862 12962 48872 13550
rect 49458 12962 49468 13550
rect 48862 12957 49468 12962
rect 48981 8285 49415 12957
rect 62648 9740 63044 9745
rect 62648 9364 62658 9740
rect 63034 9364 63044 9740
rect 62648 9359 63044 9364
rect 79162 8352 79646 8357
rect 48981 7851 50699 8285
rect 79162 7888 79172 8352
rect 79636 7888 81520 8352
rect 79162 7883 79646 7888
rect 17837 7171 20691 7605
rect 20257 -2373 20691 7171
rect 50265 -2373 50699 7851
rect 60176 1704 60544 1709
rect 60176 1382 60186 1704
rect 60534 1382 60544 1704
rect 81056 1494 81520 7888
rect 60176 1377 60544 1382
rect 60186 -294 60514 1377
rect 78734 1030 81520 1494
rect 60186 -622 62768 -294
rect 62440 -1734 62768 -622
rect 77112 -1620 77678 -1615
rect 77112 -1634 77122 -1620
rect 63096 -1734 63444 -1729
rect 62440 -2062 63106 -1734
rect 63434 -2062 63444 -1734
rect 63096 -2067 63444 -2062
rect 77094 -2058 77122 -1634
rect 77668 -1634 77678 -1620
rect 78734 -1634 79198 1030
rect 77668 -2058 79198 -1634
rect 77094 -2098 79198 -2058
rect 20257 -2807 61509 -2373
rect 17425 -8719 17879 -8714
rect 20261 -8719 20695 -2807
rect 46881 -7734 47315 -2807
rect 61075 -4119 61509 -2807
rect 61075 -4553 74008 -4119
rect 46871 -7739 47325 -7734
rect 46871 -8173 46881 -7739
rect 47315 -8173 47325 -7739
rect 46871 -8178 47325 -8173
rect 48906 -7896 49258 -7891
rect 48906 -8228 48916 -7896
rect 49248 -8228 49258 -7896
rect 48906 -8233 49258 -8228
rect 73574 -8629 74008 -4553
rect 17425 -9153 17435 -8719
rect 17869 -9153 20695 -8719
rect 73536 -8634 74018 -8629
rect 73536 -9152 73546 -8634
rect 74008 -9152 74018 -8634
rect 17425 -9158 17879 -9153
rect 73536 -9157 74018 -9152
rect -7036 -12368 -6328 -12363
rect -731 -12366 -189 -12361
rect -731 -12368 -721 -12366
rect -7036 -12898 -7026 -12368
rect -6338 -12888 -721 -12368
rect -199 -12888 -189 -12366
rect 66536 -12386 66858 -12381
rect 66536 -12404 66546 -12386
rect -6338 -12893 -189 -12888
rect 66530 -12598 66546 -12404
rect 66848 -12598 66858 -12386
rect -6338 -12898 -430 -12893
rect -7036 -12903 -6328 -12898
rect 47597 -12965 48279 -12960
rect 19335 -13021 19741 -13016
rect 19335 -13407 19345 -13021
rect 19731 -13407 19741 -13021
rect 19335 -13412 19741 -13407
rect 47597 -13627 47607 -12965
rect 48269 -13627 48279 -12965
rect 47597 -13632 48279 -13627
rect 66530 -14822 66858 -12598
rect 64424 -15150 66858 -14822
rect 17418 -16312 17766 -16307
rect 17418 -16640 17428 -16312
rect 17756 -16640 17766 -16312
rect 17418 -16645 17766 -16640
rect 48434 -16340 48782 -16335
rect 17428 -19146 17756 -16645
rect 48434 -16668 48444 -16340
rect 48772 -16668 48782 -16340
rect 48434 -16673 48782 -16668
rect 28672 -18338 29296 -18333
rect 28672 -18942 28682 -18338
rect 29286 -18942 29296 -18338
rect 28672 -18947 29296 -18942
rect 48444 -18922 48772 -16673
rect 57439 -17543 57805 -17538
rect 57439 -17889 57449 -17543
rect 57795 -17889 57805 -17543
rect 57439 -17894 57805 -17889
rect 64424 -18922 64752 -15150
rect 80404 -17382 81026 -17377
rect 80404 -18100 80414 -17382
rect 81016 -18100 81026 -17382
rect 80404 -18105 81026 -18100
rect 17428 -19474 18456 -19146
rect 48444 -19250 64752 -18922
rect 18128 -23156 18456 -19474
rect 51320 -23156 51648 -19250
rect 80316 -19874 80938 -19869
rect 80316 -20592 80326 -19874
rect 80928 -20592 80938 -19874
rect 80316 -20597 80938 -20592
rect 16792 -23438 17200 -23433
rect 16792 -23826 16802 -23438
rect 17190 -23826 17200 -23438
rect 18128 -23484 51648 -23156
rect 16792 -23831 17200 -23826
rect -7354 -24856 -6230 -24650
rect 19766 -24670 25690 -24186
rect -7354 -25568 14934 -24856
rect 19766 -24946 20250 -24670
rect 25206 -24946 25690 -24670
rect -7354 -36155 -6230 -25568
rect 14222 -28597 14934 -25568
rect 16898 -25430 20264 -24946
rect 25206 -25430 48718 -24946
rect 14174 -28602 14988 -28597
rect 14174 -29078 14184 -28602
rect 14978 -29078 14988 -28602
rect 14174 -29083 14988 -29078
rect 16898 -29661 17382 -25430
rect 48234 -29571 48718 -25430
rect 16862 -29666 17382 -29661
rect 16862 -30146 16872 -29666
rect 17352 -30146 17382 -29666
rect 48224 -29576 48728 -29571
rect 48224 -30060 48234 -29576
rect 48718 -30060 48728 -29576
rect 48224 -30065 48728 -30060
rect 16862 -30148 17382 -30146
rect 16862 -30151 17362 -30148
rect 28232 -36128 28992 -36123
rect -7380 -36160 -6206 -36155
rect -7380 -36940 -7370 -36160
rect -6216 -36940 -6206 -36160
rect 28232 -36816 28242 -36128
rect 28982 -36816 28992 -36128
rect 28232 -36821 28992 -36816
rect -7380 -36945 -6206 -36940
rect 47882 -37184 48230 -37179
rect 51320 -37184 51648 -23484
rect 62443 -27949 63157 -27944
rect 62443 -28643 62453 -27949
rect 63147 -28643 63157 -27949
rect 62443 -28648 63157 -28643
rect 55084 -31772 55706 -31767
rect 55084 -32322 55094 -31772
rect 55696 -32322 55706 -31772
rect 55084 -32327 55706 -32322
rect 47882 -37512 47892 -37184
rect 48220 -37512 51648 -37184
rect 47882 -37517 48230 -37512
<< via3 >>
rect 62658 9364 63034 9740
rect 48916 -8228 49248 -7896
rect 19345 -13407 19731 -13021
rect 47607 -13627 48269 -12965
rect 28682 -18942 29286 -18338
rect 57449 -17889 57795 -17543
rect 80414 -18100 81016 -17382
rect 80326 -20592 80928 -19874
rect 16802 -23826 17190 -23438
rect -7050 -36884 -6446 -36280
rect 28242 -36816 28982 -36128
rect 62453 -28643 63147 -27949
rect 55094 -32322 55696 -31772
<< metal4 >>
rect 62657 9740 63035 9741
rect 60396 9364 62658 9740
rect 63034 9364 63035 9740
rect 60396 5540 60772 9364
rect 62657 9363 63035 9364
rect 56628 5164 60772 5540
rect 56628 -1096 57004 5164
rect 52078 -1472 57004 -1096
rect 52078 -7880 52454 -1472
rect 48902 -7896 52454 -7880
rect 48902 -8228 48916 -7896
rect 49248 -8228 52454 -7896
rect 48902 -8256 52454 -8228
rect 47606 -12965 48270 -12964
rect 19344 -13021 19732 -13020
rect 19344 -13407 19345 -13021
rect 19731 -13407 19732 -13021
rect 19344 -13408 19732 -13407
rect 19345 -19895 19731 -13408
rect 47606 -13627 47607 -12965
rect 48269 -13627 48270 -12965
rect 47606 -13628 48270 -13627
rect 16806 -20281 19731 -19895
rect 28652 -18338 29314 -18296
rect 28652 -18942 28682 -18338
rect 29286 -18942 29314 -18338
rect 16806 -23437 17192 -20281
rect 16801 -23438 17192 -23437
rect 16801 -23826 16802 -23438
rect 17190 -23814 17192 -23438
rect 28652 -23656 29314 -18942
rect 47607 -23656 48269 -13628
rect 80413 -17382 81017 -17381
rect 80413 -17534 80414 -17382
rect 57454 -17542 80414 -17534
rect 57448 -17543 80414 -17542
rect 57448 -17889 57449 -17543
rect 57795 -17889 80414 -17543
rect 57448 -17890 80414 -17889
rect 57454 -17912 80414 -17890
rect 80413 -18100 80414 -17912
rect 81016 -18100 81017 -17382
rect 80413 -18101 81017 -18100
rect 80325 -19874 80929 -19873
rect 80325 -19944 80326 -19874
rect 69930 -20592 80326 -19944
rect 80928 -20592 80929 -19874
rect 69930 -20593 80929 -20592
rect 69930 -20596 80430 -20593
rect 69930 -20884 70582 -20596
rect 17190 -23826 17191 -23814
rect 16801 -23827 17191 -23826
rect 28652 -24318 48269 -23656
rect 62460 -21414 70582 -20884
rect 62460 -21518 76906 -21414
rect 62460 -21536 70582 -21518
rect 26917 -26711 55724 -26081
rect 26917 -29150 27547 -26711
rect 26917 -36176 27548 -29150
rect 55094 -30841 55724 -26711
rect 62460 -27948 63112 -21536
rect 70186 -21904 70290 -21536
rect 76802 -21936 76906 -21518
rect 62452 -27949 63148 -27948
rect 62452 -28643 62453 -27949
rect 63147 -28643 63148 -27949
rect 62452 -28644 63148 -28643
rect 55094 -31471 61017 -30841
rect 55094 -31771 55724 -31471
rect 55093 -31772 55724 -31771
rect 55093 -32322 55094 -31772
rect 55696 -32240 55724 -31772
rect 55696 -32322 55697 -32240
rect 55093 -32323 55697 -32322
rect 28241 -36128 28983 -36127
rect 28241 -36176 28242 -36128
rect -7051 -36280 -6445 -36279
rect -7051 -36884 -7050 -36280
rect -6446 -36884 -6445 -36280
rect 26917 -36807 28242 -36176
rect 28241 -36816 28242 -36807
rect 28982 -36816 28983 -36128
rect 28241 -36817 28983 -36816
rect -7051 -36885 -6445 -36884
rect 60387 -41107 61017 -31471
rect 66910 -40888 67014 -40726
rect 73522 -40888 73626 -40688
rect 66910 -40992 73626 -40888
rect 69804 -41107 70438 -40992
rect 60387 -41737 70439 -41107
use sky130_fd_pr__cap_mim_m3_1_L6ZKLG  sky130_fd_pr__cap_mim_m3_1_L6ZKLG_0
timestamp 1770389351
transform 1 0 70414 0 1 -31312
box -6492 -9480 6492 9480
use OFCB  x1
timestamp 1768581666
transform 1 0 958 0 1 -18688
box -914 -3502 15456 12442
use OFCB  x2
timestamp 1768581666
transform 1 0 31946 0 1 3428
box -914 -3502 15456 12442
use OFCB  x3
timestamp 1768581666
transform 1 0 31844 0 1 -18762
box -914 -3502 15456 12442
use OFCB  x4
timestamp 1768581666
transform 1 0 64098 0 1 3470
box -914 -3502 15456 12442
use OFCB  x5
timestamp 1768581666
transform 1 0 808 0 1 -39664
box -914 -3502 15456 12442
use OFCB  x6
timestamp 1768581666
transform 1 0 31770 0 1 -39668
box -914 -3502 15456 12442
use OFCB  x16
timestamp 1768581666
transform 1 0 922 0 1 3498
box -914 -3502 15456 12442
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR1
timestamp 1770460626
transform 0 1 8508 -1 0 -1089
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR2
timestamp 1770460626
transform 0 1 4324 -1 0 -22827
box -201 -1682 201 1682
use sky130_fd_pr__res_high_po_0p35_NL498X  XR3
timestamp 1770379997
transform 1 0 -2443 0 1 -6616
box -201 -642 201 642
use sky130_fd_pr__res_xhigh_po_0p35_X42PYB  XR4
timestamp 1770454287
transform 0 1 59942 -1 0 4133
box -201 -762 201 762
use sky130_fd_pr__res_xhigh_po_0p35_X42PYB  XR7
timestamp 1770454287
transform 1 0 48098 0 1 -11061
box -201 -762 201 762
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR11
timestamp 1770460626
transform 0 1 65542 -1 0 -1913
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR12
timestamp 1770460626
transform 0 1 53446 -1 0 -13789
box -201 -1682 201 1682
use sky130_fd_pr__res_high_po_0p35_NL498X  XR15
timestamp 1770379997
transform 1 0 -2441 0 1 -4862
box -201 -642 201 642
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR16
timestamp 1770460626
transform 0 1 56680 -1 0 -34077
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR17
timestamp 1770460626
transform 0 1 12576 -1 0 -1107
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR18
timestamp 1770460626
transform 0 1 4552 -1 0 -1107
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR19
timestamp 1770460626
transform 0 1 73412 -1 0 -1891
box -201 -1682 201 1682
use sky130_fd_pr__res_high_po_5p73_SWNBN6  XR20
timestamp 1770460626
transform 0 1 20344 -1 0 -38875
box -739 -852 739 852
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR21
timestamp 1770460626
transform 0 1 12936 -1 0 -22847
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR24
timestamp 1770460626
transform 0 1 8496 -1 0 -22827
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR25
timestamp 1770460626
transform 0 1 69464 -1 0 -1885
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR26
timestamp 1770460626
transform 0 1 76028 -1 0 -1041
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR27
timestamp 1770460626
transform 0 1 53432 -1 0 -15915
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR28
timestamp 1770460626
transform 0 1 53420 -1 0 -14851
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR29
timestamp 1770460626
transform 0 1 53446 -1 0 -17103
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR30
timestamp 1770460626
transform 0 1 56708 -1 0 -37021
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR32
timestamp 1770460626
transform 0 1 56680 -1 0 -35611
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_4GRPKS  XR34
timestamp 1770460626
transform 0 1 56680 -1 0 -38513
box -201 -1682 201 1682
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR35
timestamp 1770379997
transform 0 1 57384 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR36 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 58230 -1 0 -11817
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR37
timestamp 1770379997
transform 0 1 63554 -1 0 -10683
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_DBPYMX  XR38 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 63371 -1 0 -11857
box -201 -889 201 889
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR39
timestamp 1770379997
transform 0 1 67388 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR40
timestamp 1770379997
transform 0 1 68206 -1 0 -11871
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_KNJCR4  XR41
timestamp 1770379997
transform 0 1 73036 -1 0 -10689
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_MAXMKG  XR42 ~/tt10-OTA_FC/mag
timestamp 1770379997
transform 0 1 72768 -1 0 -11883
box -201 -742 201 742
<< labels >>
rlabel metal1 -3782 -33657 -3415 -5618 1 Vcm
rlabel metal1 -7774 9480 -7574 9680 1 INp
port 1 n default input
rlabel metal1 -7664 -12788 -7464 -12588 1 INm
port 2 n default input
rlabel metal1 83248 8868 83448 9068 1 OUT
port 3 n default output
rlabel metal1 83026 -17832 83226 -17632 1 Vref
port 4 n default input
rlabel metal1 83090 -25176 83290 -24976 1 ref
port 5 n default input
rlabel metal1 83116 -20314 83316 -20114 1 OUTDRL
port 6 n default output
rlabel metal1 -7558 15468 -7358 15668 1 VDD
port 7 n default bidirectional
rlabel metal1 -7710 -42968 -7510 -42768 1 GND
port 8 n default bidirectional
rlabel space 0 0 0 0 1 Vc
rlabel metal2 68300 -7601 81181 -7287 1 Vc1
rlabel metal2 74008 -9118 82585 -8732 1 Vc2
rlabel metal2 64114 -7446 64470 -5642 1 Vc
rlabel space 0 0 0 0 1 Vb
rlabel metal2 61704 -1332 61960 13166 1 Vb
<< end >>
