magic
tech sky130A
magscale 1 2
timestamp 1768572465
<< nwell >>
rect -419 -619 419 619
<< pmoslvt >>
rect -223 -400 223 400
<< pdiff >>
rect -281 388 -223 400
rect -281 -388 -269 388
rect -235 -388 -223 388
rect -281 -400 -223 -388
rect 223 388 281 400
rect 223 -388 235 388
rect 269 -388 281 388
rect 223 -400 281 -388
<< pdiffc >>
rect -269 -388 -235 388
rect 235 -388 269 388
<< nsubdiff >>
rect -383 549 -287 583
rect 287 549 383 583
rect -383 487 -349 549
rect 349 487 383 549
rect -383 -549 -349 -487
rect 349 -549 383 -487
rect -383 -583 -287 -549
rect 287 -583 383 -549
<< nsubdiffcont >>
rect -287 549 287 583
rect -383 -487 -349 487
rect 349 -487 383 487
rect -287 -583 287 -549
<< poly >>
rect -223 481 223 497
rect -223 447 -207 481
rect 207 447 223 481
rect -223 400 223 447
rect -223 -447 223 -400
rect -223 -481 -207 -447
rect 207 -481 223 -447
rect -223 -497 223 -481
<< polycont >>
rect -207 447 207 481
rect -207 -481 207 -447
<< locali >>
rect -383 549 -287 583
rect 287 549 383 583
rect -383 487 -349 549
rect 349 487 383 549
rect -223 447 -207 481
rect 207 447 223 481
rect -269 388 -235 404
rect -269 -404 -235 -388
rect 235 388 269 404
rect 235 -404 269 -388
rect -223 -481 -207 -447
rect 207 -481 223 -447
rect -383 -549 -349 -487
rect 349 -549 383 -487
rect -383 -583 -287 -549
rect 287 -583 383 -549
<< viali >>
rect -207 447 207 481
rect -269 -388 -235 388
rect 235 -388 269 388
rect -207 -481 207 -447
<< metal1 >>
rect -219 481 219 487
rect -219 447 -207 481
rect 207 447 219 481
rect -219 441 219 447
rect -275 388 -229 400
rect -275 -388 -269 388
rect -235 -388 -229 388
rect -275 -400 -229 -388
rect 229 388 275 400
rect 229 -388 235 388
rect 269 -388 275 388
rect 229 -400 275 -388
rect -219 -447 219 -441
rect -219 -481 -207 -447
rect 207 -481 219 -447
rect -219 -487 219 -481
<< properties >>
string FIXED_BBOX -366 -566 366 566
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.0 l 2.23 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
