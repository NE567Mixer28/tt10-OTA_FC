magic
tech sky130A
magscale 1 2
timestamp 1752838771
<< metal1 >>
rect 3202 16642 10312 16644
rect 3060 16636 10312 16642
rect 2708 16204 2718 16636
rect 3150 16210 10312 16636
rect 3150 16204 3160 16210
rect 3202 16208 10312 16210
rect 8698 10398 10008 10400
rect 7894 9808 7904 10398
rect 8752 9810 10008 10398
rect 30152 10232 30162 10238
rect 29564 9852 30162 10232
rect 30696 9852 30706 10238
rect 29564 9850 30698 9852
rect 8752 9808 8762 9810
rect 8438 6428 8448 7038
rect 9132 6430 11180 7038
rect 9132 6428 9142 6430
rect 4594 4258 4604 4792
rect 5134 4788 8816 4792
rect 5134 4264 10226 4788
rect 5134 4258 8816 4264
<< via1 >>
rect 2718 16204 3150 16636
rect 7904 9808 8752 10398
rect 30162 9852 30696 10238
rect 8448 6428 9132 7038
rect 4604 4258 5134 4792
<< metal2 >>
rect 2718 16636 3150 16646
rect 2718 16194 3150 16204
rect 7438 10408 8286 10410
rect 7438 10400 8752 10408
rect 8286 10398 8752 10400
rect 30162 10238 30696 10248
rect 30162 9842 30696 9852
rect 7438 9808 7904 9810
rect 7438 9800 8752 9808
rect 7904 9798 8752 9800
rect 8448 7038 9132 7048
rect 8448 6298 9132 6308
rect 4604 4792 5134 4802
rect 4604 4248 5134 4258
<< via2 >>
rect 2718 16204 3150 16636
rect 7438 10398 8286 10400
rect 7438 9810 7904 10398
rect 7904 9810 8286 10398
rect 30162 9852 30696 10238
rect 8448 6428 9132 6918
rect 8448 6308 9132 6428
rect 4604 4258 5134 4792
<< metal3 >>
rect 2708 16636 3160 16641
rect 2708 16204 2718 16636
rect 3150 16204 3160 16636
rect 2708 16199 3160 16204
rect 7428 10400 8296 10405
rect 7010 9810 7020 10400
rect 8286 9810 8296 10400
rect 30152 10238 30706 10243
rect 30152 9852 30162 10238
rect 30696 9852 30706 10238
rect 30152 9847 30706 9852
rect 7428 9805 8296 9810
rect 8438 6918 9142 6923
rect 8438 5846 8448 6918
rect 9132 5846 9142 6918
rect 4594 4792 5144 4797
rect 4594 4258 4604 4792
rect 5134 4258 5144 4792
rect 4594 4253 5144 4258
<< via3 >>
rect 2718 16204 3150 16636
rect 7020 9810 7438 10400
rect 7438 9810 7868 10400
rect 30162 9852 30696 10238
rect 8448 6308 9132 6456
rect 8448 5846 9132 6308
rect 4604 4258 5134 4792
<< metal4 >>
rect 6134 45018 6194 45152
rect 6686 45018 6746 45152
rect 7238 45018 7298 45152
rect 7790 45018 7850 45152
rect 8342 45018 8402 45152
rect 8894 45018 8954 45152
rect 9446 45018 9506 45152
rect 9998 45018 10058 45152
rect 10550 45018 10610 45152
rect 11102 45018 11162 45152
rect 11654 45018 11714 45152
rect 12206 45018 12266 45152
rect 12758 45018 12818 45152
rect 13310 45018 13370 45152
rect 13862 45018 13922 45152
rect 14414 45018 14474 45152
rect 14966 45018 15026 45152
rect 15518 45018 15578 45152
rect 16070 45018 16130 45152
rect 16622 45018 16682 45152
rect 17174 45018 17234 45152
rect 17726 45018 17786 45152
rect 18278 45018 18338 45152
rect 18830 45018 18890 45152
rect 19382 45018 19442 45152
rect 19934 45018 19994 45152
rect 20486 45018 20546 45152
rect 21038 45018 21098 45152
rect 21590 45018 21650 45152
rect 22142 45018 22202 45152
rect 22694 45018 22754 45152
rect 23246 45018 23306 45152
rect 23798 45018 23858 45152
rect 24350 45018 24410 45152
rect 24902 45018 24962 45152
rect 25454 45018 25514 45152
rect 26006 45018 26066 45152
rect 26558 45018 26618 45152
rect 27110 45018 27170 45152
rect 27662 45018 27722 45152
rect 28214 45018 28274 45152
rect 28766 45018 28826 45152
rect 29318 45018 29378 45152
rect 3710 44830 29506 45018
rect 3690 44618 29506 44830
rect 200 16634 600 44152
rect 3690 44126 4090 44618
rect 28448 44614 29506 44618
rect 3690 43982 4092 44126
rect 2717 16636 3151 16637
rect 2717 16634 2718 16636
rect 200 16204 2718 16634
rect 3150 16204 3151 16636
rect 200 16203 3151 16204
rect 200 16194 3032 16203
rect 200 1000 600 16194
rect 3692 4790 4092 43982
rect 6644 10401 7472 10404
rect 6644 10400 7869 10401
rect 6644 9810 7020 10400
rect 7868 9810 7869 10400
rect 30161 10238 30697 10239
rect 30161 9852 30162 10238
rect 30696 9852 30697 10238
rect 30161 9851 30697 9852
rect 6644 9809 7869 9810
rect 4603 4792 5135 4793
rect 4603 4790 4604 4792
rect 3692 4258 4604 4790
rect 5134 4258 5135 4792
rect 3692 974 4092 4258
rect 4603 4257 5135 4258
rect 6644 2032 7472 9809
rect 8447 6456 9133 6457
rect 8447 5992 8448 6456
rect 8438 5846 8448 5992
rect 9132 5992 9133 6456
rect 9132 5846 9162 5992
rect 8438 4038 9162 5846
rect 8444 3784 9158 4038
rect 8416 3774 26864 3784
rect 8416 2926 26910 3774
rect 6644 1966 22988 2032
rect 6644 1348 22998 1966
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22334 86 22998 1348
rect 26298 88 26910 2926
rect 30166 114 30696 9851
rect 22634 0 22814 86
rect 26498 0 26678 88
rect 30362 0 30542 114
use OFC  OFC_0
timestamp 1752750120
transform 1 0 6786 0 1 4062
box 2996 206 22976 12566
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 3692 974 4092 44126 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
