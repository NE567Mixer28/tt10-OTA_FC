magic
tech sky130A
magscale 1 2
timestamp 1770460626
<< pwell >>
rect -739 -852 739 852
<< psubdiff >>
rect -703 782 -607 816
rect 607 782 703 816
rect -703 720 -669 782
rect 669 720 703 782
rect -703 -782 -669 -720
rect 669 -782 703 -720
rect -703 -816 -607 -782
rect 607 -816 703 -782
<< psubdiffcont >>
rect -607 782 607 816
rect -703 -720 -669 720
rect 669 -720 703 720
rect -607 -816 607 -782
<< xpolycontact >>
rect -573 254 573 686
rect -573 -686 573 -254
<< ppolyres >>
rect -573 -254 573 254
<< locali >>
rect -703 782 -607 816
rect 607 782 703 816
rect -703 720 -669 782
rect 669 720 703 782
rect -703 -782 -669 -720
rect 669 -782 703 -720
rect -703 -816 -607 -782
rect 607 -816 703 -782
<< viali >>
rect -557 271 557 668
rect -557 -668 557 -271
<< metal1 >>
rect -569 668 569 674
rect -569 271 -557 668
rect 557 271 569 668
rect -569 265 569 271
rect -569 -271 569 -265
rect -569 -668 -557 -271
rect 557 -668 569 -271
rect -569 -674 569 -668
<< properties >>
string FIXED_BBOX -686 -799 686 799
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 5.730 l 2.7 m 1 nx 1 wmin 5.730 lmin 0.50 rho 319.8 val 218.691 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
