** sch_path: /home/ttuser/tt10-OTA_FC/xschem/ecg.sch
.subckt ecg VDD GND INp INm Odrl OUT ref
*.PININFO VDD:B GND:B INp:I INm:I Odrl:O OUT:O ref:I
XR3 Vcm net3 GND sky130_fd_pr__res_high_po_0p35 L=0.4 mult=1 m=1
XR15 Vcm net4 GND sky130_fd_pr__res_high_po_0p35 L=0.4 mult=1 m=1
XR18 net3 net7 GND sky130_fd_pr__res_xhigh_po_0p35 L=10 mult=1 m=1
XR20 net6 net5 GND sky130_fd_pr__res_high_po_5p73 L=2.7 mult=1 m=1
XR17 net8 out1 GND sky130_fd_pr__res_xhigh_po_0p35 L=6.2 mult=1 m=1
XR1 net7 net8 GND sky130_fd_pr__res_xhigh_po_0p35 L=10 mult=1 m=1
XR2 net4 net9 GND sky130_fd_pr__res_xhigh_po_0p35 L=10 mult=1 m=1
XR21 net10 out2 GND sky130_fd_pr__res_xhigh_po_0p35 L=6.2 mult=1 m=1
XR24 net9 net10 GND sky130_fd_pr__res_xhigh_po_0p35 L=10 mult=1 m=1
XR4 out12 net2 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.8 mult=1 m=1
XR7 out22 net1 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.8 mult=1 m=1
XR11 net2 net11 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR19 net12 net13 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR25 net11 net12 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR26 net13 OUT GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR12 net1 net14 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR27 net15 net16 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR28 net14 net15 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR29 net16 ref GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR16 net5 net17 GND sky130_fd_pr__res_xhigh_po_0p35 L=8.7 mult=1 m=1
XR30 net17 Odrl GND sky130_fd_pr__res_xhigh_po_0p35 L=8.7 mult=1 m=1
XC2 net5 Odrl sky130_fd_pr__cap_mim_m3_1 W=71 L=71 m=1
x1 VDD GND out1 net3 INp OFC
x2 VDD GND out2 net4 INm OFC
x3 VDD GND out12 out12 out1 OFC
x4 VDD GND out22 out22 out2 OFC
x5 VDD GND OUT net2 net1 OFC
x6 VDD GND net6 net6 Vcm OFC
x7 VDD GND Odrl net5 ref OFC
.ends

* expanding   symbol:  OFC.sym # of pins=5
** sym_path: /home/ttuser/tt10-OTA_FC/xschem/OFC.sym
** sch_path: /home/ttuser/tt10-OTA_FC/xschem/OFC.sch
.subckt OFC VDD VSS OUT INm INp
*.PININFO VDD:B VSS:B INp:I INm:I OUT:O
XM11 S Vb VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=60 nf=6 m=2
XM1 D1 INp S S sky130_fd_pr__pfet_01v8_lvt L=10 W=25 nf=2 m=2
XM2 D2 INm S S sky130_fd_pr__pfet_01v8_lvt L=10 W=25 nf=2 m=2
XM3 OUT Vc1 D2 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM4 D2 Vc VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2.8 nf=1 m=1
XM5 D1 Vc VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2.8 nf=1 m=1
XM6 G Vc1 D1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 m=1
XM7 G Vc2 D9 D9 sky130_fd_pr__pfet_01v8_lvt L=2.23 W=3 nf=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2.23 W=4 nf=1 m=1
XM8 D10 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2.23 W=4 nf=1 m=1
XM10 OUT Vc2 D10 D10 sky130_fd_pr__pfet_01v8_lvt L=2.23 W=3 nf=1 m=1
XR2 Vb VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR3 VSS Vb VSS sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR1 Vc VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR4 VSS Vc VSS sky130_fd_pr__res_xhigh_po_0p35 L=3.07 mult=1 m=1
XR5 Vc1 VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR6 VSS Vc1 VSS sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR7 Vc2 VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR8 VSS Vc2 VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.6 mult=1 m=1
.ends

.end
