magic
tech sky130A
magscale 1 2
timestamp 1768572465
<< nwell >>
rect -941 -2337 941 2337
<< pmoslvt >>
rect -745 118 -545 2118
rect -487 118 -287 2118
rect -229 118 -29 2118
rect 29 118 229 2118
rect 287 118 487 2118
rect 545 118 745 2118
rect -745 -2118 -545 -118
rect -487 -2118 -287 -118
rect -229 -2118 -29 -118
rect 29 -2118 229 -118
rect 287 -2118 487 -118
rect 545 -2118 745 -118
<< pdiff >>
rect -803 2106 -745 2118
rect -803 130 -791 2106
rect -757 130 -745 2106
rect -803 118 -745 130
rect -545 2106 -487 2118
rect -545 130 -533 2106
rect -499 130 -487 2106
rect -545 118 -487 130
rect -287 2106 -229 2118
rect -287 130 -275 2106
rect -241 130 -229 2106
rect -287 118 -229 130
rect -29 2106 29 2118
rect -29 130 -17 2106
rect 17 130 29 2106
rect -29 118 29 130
rect 229 2106 287 2118
rect 229 130 241 2106
rect 275 130 287 2106
rect 229 118 287 130
rect 487 2106 545 2118
rect 487 130 499 2106
rect 533 130 545 2106
rect 487 118 545 130
rect 745 2106 803 2118
rect 745 130 757 2106
rect 791 130 803 2106
rect 745 118 803 130
rect -803 -130 -745 -118
rect -803 -2106 -791 -130
rect -757 -2106 -745 -130
rect -803 -2118 -745 -2106
rect -545 -130 -487 -118
rect -545 -2106 -533 -130
rect -499 -2106 -487 -130
rect -545 -2118 -487 -2106
rect -287 -130 -229 -118
rect -287 -2106 -275 -130
rect -241 -2106 -229 -130
rect -287 -2118 -229 -2106
rect -29 -130 29 -118
rect -29 -2106 -17 -130
rect 17 -2106 29 -130
rect -29 -2118 29 -2106
rect 229 -130 287 -118
rect 229 -2106 241 -130
rect 275 -2106 287 -130
rect 229 -2118 287 -2106
rect 487 -130 545 -118
rect 487 -2106 499 -130
rect 533 -2106 545 -130
rect 487 -2118 545 -2106
rect 745 -130 803 -118
rect 745 -2106 757 -130
rect 791 -2106 803 -130
rect 745 -2118 803 -2106
<< pdiffc >>
rect -791 130 -757 2106
rect -533 130 -499 2106
rect -275 130 -241 2106
rect -17 130 17 2106
rect 241 130 275 2106
rect 499 130 533 2106
rect 757 130 791 2106
rect -791 -2106 -757 -130
rect -533 -2106 -499 -130
rect -275 -2106 -241 -130
rect -17 -2106 17 -130
rect 241 -2106 275 -130
rect 499 -2106 533 -130
rect 757 -2106 791 -130
<< nsubdiff >>
rect -905 2267 -809 2301
rect 809 2267 905 2301
rect -905 2205 -871 2267
rect 871 2205 905 2267
rect -905 -2267 -871 -2205
rect 871 -2267 905 -2205
rect -905 -2301 -809 -2267
rect 809 -2301 905 -2267
<< nsubdiffcont >>
rect -809 2267 809 2301
rect -905 -2205 -871 2205
rect 871 -2205 905 2205
rect -809 -2301 809 -2267
<< poly >>
rect -745 2199 -545 2215
rect -745 2165 -729 2199
rect -561 2165 -545 2199
rect -745 2118 -545 2165
rect -487 2199 -287 2215
rect -487 2165 -471 2199
rect -303 2165 -287 2199
rect -487 2118 -287 2165
rect -229 2199 -29 2215
rect -229 2165 -213 2199
rect -45 2165 -29 2199
rect -229 2118 -29 2165
rect 29 2199 229 2215
rect 29 2165 45 2199
rect 213 2165 229 2199
rect 29 2118 229 2165
rect 287 2199 487 2215
rect 287 2165 303 2199
rect 471 2165 487 2199
rect 287 2118 487 2165
rect 545 2199 745 2215
rect 545 2165 561 2199
rect 729 2165 745 2199
rect 545 2118 745 2165
rect -745 71 -545 118
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 118
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -118 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -118 745 -71
rect -745 -2165 -545 -2118
rect -745 -2199 -729 -2165
rect -561 -2199 -545 -2165
rect -745 -2215 -545 -2199
rect -487 -2165 -287 -2118
rect -487 -2199 -471 -2165
rect -303 -2199 -287 -2165
rect -487 -2215 -287 -2199
rect -229 -2165 -29 -2118
rect -229 -2199 -213 -2165
rect -45 -2199 -29 -2165
rect -229 -2215 -29 -2199
rect 29 -2165 229 -2118
rect 29 -2199 45 -2165
rect 213 -2199 229 -2165
rect 29 -2215 229 -2199
rect 287 -2165 487 -2118
rect 287 -2199 303 -2165
rect 471 -2199 487 -2165
rect 287 -2215 487 -2199
rect 545 -2165 745 -2118
rect 545 -2199 561 -2165
rect 729 -2199 745 -2165
rect 545 -2215 745 -2199
<< polycont >>
rect -729 2165 -561 2199
rect -471 2165 -303 2199
rect -213 2165 -45 2199
rect 45 2165 213 2199
rect 303 2165 471 2199
rect 561 2165 729 2199
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect -729 -2199 -561 -2165
rect -471 -2199 -303 -2165
rect -213 -2199 -45 -2165
rect 45 -2199 213 -2165
rect 303 -2199 471 -2165
rect 561 -2199 729 -2165
<< locali >>
rect -905 2267 -809 2301
rect 809 2267 905 2301
rect -905 2205 -871 2267
rect 871 2205 905 2267
rect -745 2165 -729 2199
rect -561 2165 -545 2199
rect -487 2165 -471 2199
rect -303 2165 -287 2199
rect -229 2165 -213 2199
rect -45 2165 -29 2199
rect 29 2165 45 2199
rect 213 2165 229 2199
rect 287 2165 303 2199
rect 471 2165 487 2199
rect 545 2165 561 2199
rect 729 2165 745 2199
rect -791 2106 -757 2122
rect -791 114 -757 130
rect -533 2106 -499 2122
rect -533 114 -499 130
rect -275 2106 -241 2122
rect -275 114 -241 130
rect -17 2106 17 2122
rect -17 114 17 130
rect 241 2106 275 2122
rect 241 114 275 130
rect 499 2106 533 2122
rect 499 114 533 130
rect 757 2106 791 2122
rect 757 114 791 130
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect -791 -130 -757 -114
rect -791 -2122 -757 -2106
rect -533 -130 -499 -114
rect -533 -2122 -499 -2106
rect -275 -130 -241 -114
rect -275 -2122 -241 -2106
rect -17 -130 17 -114
rect -17 -2122 17 -2106
rect 241 -130 275 -114
rect 241 -2122 275 -2106
rect 499 -130 533 -114
rect 499 -2122 533 -2106
rect 757 -130 791 -114
rect 757 -2122 791 -2106
rect -745 -2199 -729 -2165
rect -561 -2199 -545 -2165
rect -487 -2199 -471 -2165
rect -303 -2199 -287 -2165
rect -229 -2199 -213 -2165
rect -45 -2199 -29 -2165
rect 29 -2199 45 -2165
rect 213 -2199 229 -2165
rect 287 -2199 303 -2165
rect 471 -2199 487 -2165
rect 545 -2199 561 -2165
rect 729 -2199 745 -2165
rect -905 -2267 -871 -2205
rect 871 -2267 905 -2205
rect -905 -2301 -809 -2267
rect 809 -2301 905 -2267
<< viali >>
rect -729 2165 -561 2199
rect -471 2165 -303 2199
rect -213 2165 -45 2199
rect 45 2165 213 2199
rect 303 2165 471 2199
rect 561 2165 729 2199
rect -791 130 -757 2106
rect -533 130 -499 2106
rect -275 130 -241 2106
rect -17 130 17 2106
rect 241 130 275 2106
rect 499 130 533 2106
rect 757 130 791 2106
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect -791 -2106 -757 -130
rect -533 -2106 -499 -130
rect -275 -2106 -241 -130
rect -17 -2106 17 -130
rect 241 -2106 275 -130
rect 499 -2106 533 -130
rect 757 -2106 791 -130
rect -729 -2199 -561 -2165
rect -471 -2199 -303 -2165
rect -213 -2199 -45 -2165
rect 45 -2199 213 -2165
rect 303 -2199 471 -2165
rect 561 -2199 729 -2165
<< metal1 >>
rect -741 2199 -549 2205
rect -741 2165 -729 2199
rect -561 2165 -549 2199
rect -741 2159 -549 2165
rect -483 2199 -291 2205
rect -483 2165 -471 2199
rect -303 2165 -291 2199
rect -483 2159 -291 2165
rect -225 2199 -33 2205
rect -225 2165 -213 2199
rect -45 2165 -33 2199
rect -225 2159 -33 2165
rect 33 2199 225 2205
rect 33 2165 45 2199
rect 213 2165 225 2199
rect 33 2159 225 2165
rect 291 2199 483 2205
rect 291 2165 303 2199
rect 471 2165 483 2199
rect 291 2159 483 2165
rect 549 2199 741 2205
rect 549 2165 561 2199
rect 729 2165 741 2199
rect 549 2159 741 2165
rect -797 2106 -751 2118
rect -797 130 -791 2106
rect -757 130 -751 2106
rect -797 118 -751 130
rect -539 2106 -493 2118
rect -539 130 -533 2106
rect -499 130 -493 2106
rect -539 118 -493 130
rect -281 2106 -235 2118
rect -281 130 -275 2106
rect -241 130 -235 2106
rect -281 118 -235 130
rect -23 2106 23 2118
rect -23 130 -17 2106
rect 17 130 23 2106
rect -23 118 23 130
rect 235 2106 281 2118
rect 235 130 241 2106
rect 275 130 281 2106
rect 235 118 281 130
rect 493 2106 539 2118
rect 493 130 499 2106
rect 533 130 539 2106
rect 493 118 539 130
rect 751 2106 797 2118
rect 751 130 757 2106
rect 791 130 797 2106
rect 751 118 797 130
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect -797 -130 -751 -118
rect -797 -2106 -791 -130
rect -757 -2106 -751 -130
rect -797 -2118 -751 -2106
rect -539 -130 -493 -118
rect -539 -2106 -533 -130
rect -499 -2106 -493 -130
rect -539 -2118 -493 -2106
rect -281 -130 -235 -118
rect -281 -2106 -275 -130
rect -241 -2106 -235 -130
rect -281 -2118 -235 -2106
rect -23 -130 23 -118
rect -23 -2106 -17 -130
rect 17 -2106 23 -130
rect -23 -2118 23 -2106
rect 235 -130 281 -118
rect 235 -2106 241 -130
rect 275 -2106 281 -130
rect 235 -2118 281 -2106
rect 493 -130 539 -118
rect 493 -2106 499 -130
rect 533 -2106 539 -130
rect 493 -2118 539 -2106
rect 751 -130 797 -118
rect 751 -2106 757 -130
rect 791 -2106 797 -130
rect 751 -2118 797 -2106
rect -741 -2165 -549 -2159
rect -741 -2199 -729 -2165
rect -561 -2199 -549 -2165
rect -741 -2205 -549 -2199
rect -483 -2165 -291 -2159
rect -483 -2199 -471 -2165
rect -303 -2199 -291 -2165
rect -483 -2205 -291 -2199
rect -225 -2165 -33 -2159
rect -225 -2199 -213 -2165
rect -45 -2199 -33 -2165
rect -225 -2205 -33 -2199
rect 33 -2165 225 -2159
rect 33 -2199 45 -2165
rect 213 -2199 225 -2165
rect 33 -2205 225 -2199
rect 291 -2165 483 -2159
rect 291 -2199 303 -2165
rect 471 -2199 483 -2165
rect 291 -2205 483 -2199
rect 549 -2165 741 -2159
rect 549 -2199 561 -2165
rect 729 -2199 741 -2165
rect 549 -2205 741 -2199
<< properties >>
string FIXED_BBOX -888 -2284 888 2284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
