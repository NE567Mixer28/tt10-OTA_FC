magic
tech sky130A
magscale 1 2
timestamp 1770379997
<< pwell >>
rect -201 -889 201 889
<< psubdiff >>
rect -165 819 -69 853
rect 69 819 165 853
rect -165 757 -131 819
rect 131 757 165 819
rect -165 -819 -131 -757
rect 131 -819 165 -757
rect -165 -853 -69 -819
rect 69 -853 165 -819
<< psubdiffcont >>
rect -69 819 69 853
rect -165 -757 -131 757
rect 131 -757 165 757
rect -69 -853 69 -819
<< xpolycontact >>
rect -35 291 35 723
rect -35 -723 35 -291
<< xpolyres >>
rect -35 -291 35 291
<< locali >>
rect -165 819 -69 853
rect 69 819 165 853
rect -165 757 -131 819
rect 131 757 165 819
rect -165 -819 -131 -757
rect 131 -819 165 -757
rect -165 -853 -69 -819
rect 69 -853 165 -819
<< viali >>
rect -19 308 19 705
rect -19 -705 19 -308
<< metal1 >>
rect -25 705 25 717
rect -25 308 -19 705
rect 19 308 25 705
rect -25 296 25 308
rect -25 -308 25 -296
rect -25 -705 -19 -308
rect 19 -705 25 -308
rect -25 -717 25 -705
<< properties >>
string FIXED_BBOX -148 -836 148 836
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.07 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 18.618k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
