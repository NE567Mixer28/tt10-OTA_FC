magic
tech sky130A
magscale 1 2
timestamp 1770460626
<< pwell >>
rect -201 -1682 201 1682
<< psubdiff >>
rect -165 1612 -69 1646
rect 69 1612 165 1646
rect -165 1550 -131 1612
rect 131 1550 165 1612
rect -165 -1612 -131 -1550
rect 131 -1612 165 -1550
rect -165 -1646 -69 -1612
rect 69 -1646 165 -1612
<< psubdiffcont >>
rect -69 1612 69 1646
rect -165 -1550 -131 1550
rect 131 -1550 165 1550
rect -69 -1646 69 -1612
<< xpolycontact >>
rect -35 1084 35 1516
rect -35 -1516 35 -1084
<< xpolyres >>
rect -35 -1084 35 1084
<< locali >>
rect -165 1612 -69 1646
rect 69 1612 165 1646
rect -165 1550 -131 1612
rect 131 1550 165 1612
rect -165 -1612 -131 -1550
rect 131 -1612 165 -1550
rect -165 -1646 -69 -1612
rect 69 -1646 165 -1612
<< viali >>
rect -19 1101 19 1498
rect -19 -1498 19 -1101
<< metal1 >>
rect -25 1498 25 1510
rect -25 1101 -19 1498
rect 19 1101 25 1498
rect -25 1089 25 1101
rect -25 -1101 25 -1089
rect -25 -1498 -19 -1101
rect 19 -1498 25 -1101
rect -25 -1510 25 -1498
<< properties >>
string FIXED_BBOX -148 -1629 148 1629
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 11 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 63.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
