magic
tech sky130A
magscale 1 2
timestamp 1768572465
<< nwell >>
rect -419 -604 419 604
<< pmoslvt >>
rect -223 -385 223 385
<< pdiff >>
rect -281 373 -223 385
rect -281 -373 -269 373
rect -235 -373 -223 373
rect -281 -385 -223 -373
rect 223 373 281 385
rect 223 -373 235 373
rect 269 -373 281 373
rect 223 -385 281 -373
<< pdiffc >>
rect -269 -373 -235 373
rect 235 -373 269 373
<< nsubdiff >>
rect -383 534 -287 568
rect 287 534 383 568
rect -383 472 -349 534
rect 349 472 383 534
rect -383 -534 -349 -472
rect 349 -534 383 -472
rect -383 -568 -287 -534
rect 287 -568 383 -534
<< nsubdiffcont >>
rect -287 534 287 568
rect -383 -472 -349 472
rect 349 -472 383 472
rect -287 -568 287 -534
<< poly >>
rect -223 466 223 482
rect -223 432 -207 466
rect 207 432 223 466
rect -223 385 223 432
rect -223 -432 223 -385
rect -223 -466 -207 -432
rect 207 -466 223 -432
rect -223 -482 223 -466
<< polycont >>
rect -207 432 207 466
rect -207 -466 207 -432
<< locali >>
rect -383 534 -287 568
rect 287 534 383 568
rect -383 472 -349 534
rect 349 472 383 534
rect -223 432 -207 466
rect 207 432 223 466
rect -269 373 -235 389
rect -269 -389 -235 -373
rect 235 373 269 389
rect 235 -389 269 -373
rect -223 -466 -207 -432
rect 207 -466 223 -432
rect -383 -534 -349 -472
rect 349 -534 383 -472
rect -383 -568 -287 -534
rect 287 -568 383 -534
<< viali >>
rect -207 432 207 466
rect -269 -373 -235 373
rect 235 -373 269 373
rect -207 -466 207 -432
<< metal1 >>
rect -219 466 219 472
rect -219 432 -207 466
rect 207 432 219 466
rect -219 426 219 432
rect -275 373 -229 385
rect -275 -373 -269 373
rect -235 -373 -229 373
rect -275 -385 -229 -373
rect 229 373 275 385
rect 229 -373 235 373
rect 269 -373 275 373
rect 229 -385 275 -373
rect -219 -432 219 -426
rect -219 -466 -207 -432
rect 207 -466 219 -432
rect -219 -472 219 -466
<< properties >>
string FIXED_BBOX -366 -551 366 551
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 3.85 l 2.23 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
