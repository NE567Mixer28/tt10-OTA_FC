magic
tech sky130A
magscale 1 2
timestamp 1770379997
<< error_p >>
rect -35 34 35 36
<< pwell >>
rect -201 -632 201 632
<< psubdiff >>
rect -165 562 -69 596
rect 69 562 165 596
rect -165 500 -131 562
rect 131 500 165 562
rect -165 -562 -131 -500
rect 131 -562 165 -500
rect -165 -596 -69 -562
rect 69 -596 165 -562
<< psubdiffcont >>
rect -69 562 69 596
rect -165 -500 -131 500
rect 131 -500 165 500
rect -69 -596 69 -562
<< xpolycontact >>
rect -35 34 35 466
rect -35 -466 35 -34
<< ppolyres >>
rect -35 -34 35 34
<< locali >>
rect -165 562 -69 596
rect 69 562 165 596
rect -165 500 -131 562
rect 131 500 165 562
rect -165 -562 -131 -500
rect 131 -562 165 -500
rect -165 -596 -69 -562
rect 69 -596 165 -562
<< viali >>
rect -19 51 19 448
rect -19 -448 19 -51
<< metal1 >>
rect -25 448 25 460
rect -25 51 -19 448
rect 19 51 25 448
rect -25 39 25 51
rect -25 -51 25 -39
rect -25 -448 -19 -51
rect 19 -448 25 -51
rect -25 -460 25 -448
<< properties >>
string FIXED_BBOX -148 -579 148 579
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.50 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 1.57k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
