** sch_path: /home/ttuser/tt10-OTA_FC/xschem/ecg.sch
.subckt ecg INp INm OUT Vref OUTDRL ref VDD GND
*.PININFO INp:I INm:I OUT:O Vref:I OUTDRL:O ref:I VDD:B GND:B
XR3 Vcm net3 GND sky130_fd_pr__res_high_po_0p35 L=0.6 mult=1 m=1
XR15 Vcm net4 GND sky130_fd_pr__res_high_po_0p35 L=0.6 mult=1 m=1
XR18 net3 net7 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR20 net6 net5 GND sky130_fd_pr__res_high_po_5p73 L=2.7 mult=1 m=1
XR17 net8 out1 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR1 net7 net8 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR2 net4 net9 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR21 net10 out2 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR24 net9 net10 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR4 out12 net2 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.8 mult=1 m=1
XR7 out22 net1 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.8 mult=1 m=1
XR11 net2 net11 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR19 net12 net13 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR25 net11 net12 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR26 net13 OUT GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR12 net1 net14 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR27 net15 net16 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR28 net14 net15 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR29 net16 Vref GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XC2 net5 OUTDRL sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=6 m=6
XR16 net5 net17 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR30 net18 net19 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR32 net17 net18 GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
XR34 net19 OUTDRL GND sky130_fd_pr__res_xhigh_po_0p35 L=11 mult=1 m=1
x16 Vb VDD GND Vc2 out1 INp net3 Vc1 Vc OFCB
x1 Vb VDD GND Vc2 out2 INm net4 Vc1 Vc OFCB
x2 Vb VDD GND Vc2 out12 out1 out12 Vc1 Vc OFCB
x3 Vb VDD GND Vc2 out22 out2 out22 Vc1 Vc OFCB
x4 Vb VDD GND Vc2 OUT net1 net2 Vc1 Vc OFCB
x5 Vb VDD GND Vc2 net6 Vcm net6 Vc1 Vc OFCB
x6 Vb VDD GND Vc2 OUTDRL ref net5 Vc1 Vc OFCB
XR35 Vb VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR36 GND Vb GND sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR37 Vc VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR38 GND Vc GND sky130_fd_pr__res_xhigh_po_0p35 L=3.07 mult=1 m=1
XR39 Vc1 VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR40 GND Vc1 GND sky130_fd_pr__res_xhigh_po_0p35 L=13.2 mult=1 m=1
XR41 Vc2 VDD GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR42 GND Vc2 GND sky130_fd_pr__res_xhigh_po_0p35 L=1.6 mult=1 m=1
.ends

* expanding   symbol:  OFCB.sym # of pins=9
** sym_path: /home/ttuser/tt10-OTA_FC/xschem/OFCB.sym
** sch_path: /home/ttuser/tt10-OTA_FC/xschem/OFCB.sch
.subckt OFCB Vb VDD GND Vc2 OUT INp INm Vc1 Vc
*.PININFO VDD:B GND:B OUT:O INp:I INm:I Vc2:B Vc1:B Vc:B Vb:B
XM11 S Vb VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=60 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM1 D1 INp S S sky130_fd_pr__pfet_01v8_lvt L=10 W=25 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 D2 INm S S sky130_fd_pr__pfet_01v8_lvt L=10 W=25 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 OUT Vc1 D2 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 D2 Vc GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=2.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 D1 Vc GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=2.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 G Vc1 D1 GND sky130_fd_pr__nfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 G Vc2 D9 D9 sky130_fd_pr__pfet_01v8_lvt L=2.23 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 D9 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2.23 W=3.85 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 D10 G VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2.23 W=3.85 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT Vc2 D10 D10 sky130_fd_pr__pfet_01v8_lvt L=2.23 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 OUT D1 sky130_fd_pr__cap_mim_m3_1 W=22.4 L=22.4 MF=2 m=2
.ends

.end
