magic
tech sky130A
magscale 1 2
timestamp 1753192428
<< viali >>
rect 15134 11772 15338 11840
rect 17012 11764 17218 11830
rect 8350 11482 8616 11574
rect 12102 11568 12190 11716
rect 21428 11430 21504 11538
rect 20186 11304 20346 11362
rect 13730 10900 13820 10986
rect 22110 10962 22192 11112
rect 20186 10820 20346 10912
rect 15106 10614 15344 10684
rect 16990 10606 17232 10678
rect 21736 10438 21854 10516
rect 7656 8178 7808 8242
rect 15496 8146 15722 8214
rect 21738 6746 21854 6806
rect 21734 2732 21818 2802
rect 13978 2496 14102 2538
rect 18110 2102 18214 2170
rect 13970 1620 14066 1672
rect 18106 1634 18212 1694
rect 13568 1126 13814 1182
rect 17752 1146 17938 1214
rect 21060 1042 21174 1116
rect 21714 1050 21830 1124
<< metal1 >>
rect 11972 12564 20358 12566
rect 11972 12562 22964 12564
rect 3240 12150 22964 12562
rect 5944 12068 7200 12150
rect 5936 11698 5946 12068
rect 7362 11698 7372 12068
rect 8236 11574 8788 12150
rect 10230 11612 10600 12150
rect 11972 12138 22964 12150
rect 15006 11840 15470 12138
rect 15006 11772 15134 11840
rect 15338 11772 15470 11840
rect 12096 11716 12196 11728
rect 12328 11716 13630 11718
rect 8236 11536 8350 11574
rect 8338 11482 8350 11536
rect 8616 11536 8788 11574
rect 8616 11482 8628 11536
rect 8338 11476 8628 11482
rect 5236 11342 5246 11454
rect 5628 11342 5638 11454
rect 6468 11102 6478 11214
rect 6860 11102 6870 11214
rect 5228 10850 5238 10954
rect 5636 10850 5646 10954
rect 6472 10596 6482 10708
rect 6864 10596 6874 10708
rect 5224 10334 5234 10424
rect 5636 10334 5646 10424
rect 6478 10080 6488 10192
rect 6870 10080 6880 10192
rect 7222 9910 7358 11368
rect 7630 11354 7640 11466
rect 8022 11354 8032 11466
rect 11652 11412 11962 11668
rect 12096 11568 12102 11716
rect 12190 11568 13630 11716
rect 15006 11686 15470 11772
rect 16894 11830 17358 12138
rect 20094 12118 22964 12138
rect 16894 11764 17012 11830
rect 17218 11764 17358 11830
rect 16894 11680 17358 11764
rect 12096 11556 13630 11568
rect 12112 11554 13630 11556
rect 10230 11350 12040 11412
rect 9722 11346 9872 11350
rect 9460 11308 9872 11346
rect 10228 11308 12040 11350
rect 9460 11260 12040 11308
rect 12328 11280 13630 11554
rect 15700 11572 16650 11606
rect 15700 11346 16012 11572
rect 16350 11346 16650 11572
rect 15700 11282 16650 11346
rect 9460 11210 10600 11260
rect 8804 11088 8814 11200
rect 9196 11088 9206 11200
rect 9722 11166 10600 11210
rect 9722 11138 9872 11166
rect 9722 11096 9868 11138
rect 9470 10960 9868 11096
rect 7630 10840 7640 10952
rect 8022 10840 8032 10952
rect 9722 10844 9868 10960
rect 10228 10922 10600 11166
rect 13300 10992 13624 11280
rect 19584 11234 19922 11502
rect 20982 11476 21292 12118
rect 21422 11546 21510 11550
rect 21418 11544 21892 11546
rect 21418 11538 22018 11544
rect 20178 11368 20366 11370
rect 20174 11362 20366 11368
rect 20174 11304 20186 11362
rect 20346 11304 20366 11362
rect 20174 11298 20366 11304
rect 18284 11232 19922 11234
rect 13298 10988 13624 10992
rect 13718 10988 13832 10992
rect 13298 10986 13836 10988
rect 13298 10960 13730 10986
rect 9462 10708 9868 10844
rect 8804 10580 8814 10692
rect 9196 10580 9206 10692
rect 9722 10570 9868 10708
rect 13296 10900 13730 10960
rect 13820 10900 13836 10986
rect 13296 10898 13836 10900
rect 13296 10622 13622 10898
rect 13718 10894 13832 10898
rect 7630 10328 7640 10440
rect 8022 10328 8032 10440
rect 9470 10434 9868 10570
rect 9722 10320 9868 10434
rect 13290 10540 13622 10622
rect 15016 10684 15466 11196
rect 15016 10614 15106 10684
rect 15344 10614 15466 10684
rect 13290 10350 13616 10540
rect 15016 10522 15466 10614
rect 16932 10678 17318 11188
rect 16932 10606 16990 10678
rect 17232 10606 17318 10678
rect 16932 10506 17318 10606
rect 18078 11040 19922 11232
rect 9466 10184 9868 10320
rect 8804 10066 8814 10178
rect 9196 10066 9206 10178
rect 9722 10056 9868 10184
rect 5216 9828 5226 9894
rect 5636 9828 5646 9894
rect 7630 9814 7640 9926
rect 8022 9814 8032 9926
rect 9462 9920 9868 10056
rect 12202 10024 12212 10350
rect 12602 10036 13616 10350
rect 15598 10118 16754 10436
rect 18078 10430 19218 11040
rect 19584 10694 19922 11040
rect 20178 11178 20366 11298
rect 21030 11200 21268 11476
rect 21418 11430 21428 11538
rect 21504 11430 22018 11538
rect 22216 11432 22412 12118
rect 21418 11422 22018 11430
rect 21422 11418 21510 11422
rect 20178 10918 20662 11178
rect 20174 10912 20662 10918
rect 20174 10820 20186 10912
rect 20346 10820 20662 10912
rect 20174 10814 20662 10820
rect 20314 10682 20662 10814
rect 17468 10116 19218 10430
rect 18078 10112 19218 10116
rect 18078 10110 18418 10112
rect 12602 10024 13610 10036
rect 15008 9736 15378 10020
rect 7550 9526 8072 9530
rect 7540 9306 7550 9526
rect 8068 9306 8078 9526
rect 7550 8998 8072 9306
rect 11404 9290 11414 9704
rect 11702 9698 11990 9704
rect 15008 9698 16012 9736
rect 11702 9496 16012 9698
rect 16354 9496 16364 9736
rect 16872 9732 17346 10030
rect 21030 9854 21420 11200
rect 21628 11112 22018 11422
rect 22104 11112 22198 11124
rect 21628 10962 22110 11112
rect 22192 10962 22202 11112
rect 21628 10944 22202 10962
rect 21628 10548 22018 10944
rect 21716 10516 21896 10548
rect 21716 10442 21736 10516
rect 21724 10438 21736 10442
rect 21854 10442 21896 10516
rect 21854 10438 21866 10442
rect 21724 10432 21866 10438
rect 21742 10002 21752 10288
rect 21852 10020 22312 10288
rect 21852 10002 21862 10020
rect 16870 9718 18746 9732
rect 11702 9482 16354 9496
rect 11702 9352 15332 9482
rect 11702 9290 11712 9352
rect 11904 9346 15332 9352
rect 16870 9356 20510 9718
rect 21024 9684 21034 9854
rect 21190 9740 21420 9854
rect 21190 9722 21268 9740
rect 21190 9684 21200 9722
rect 16870 9346 18746 9356
rect 5488 8994 10862 8998
rect 11256 8996 11412 8998
rect 11256 8994 14380 8996
rect 17552 8994 19296 9004
rect 5488 8984 19296 8994
rect 5488 8626 10382 8984
rect 10854 8976 19296 8984
rect 10854 8626 19324 8976
rect 5488 8554 19324 8626
rect 5488 8534 11412 8554
rect 5488 8530 11308 8534
rect 5488 8430 10862 8530
rect 13398 8448 19324 8554
rect 5532 8072 7262 8430
rect 7664 8248 7808 8430
rect 7644 8242 7820 8248
rect 7644 8178 7656 8242
rect 7808 8178 7820 8242
rect 7644 8172 7820 8178
rect 8266 8090 9996 8430
rect 13398 8052 15128 8448
rect 15494 8220 15724 8448
rect 16138 8430 19324 8448
rect 15484 8214 15734 8220
rect 15484 8146 15496 8214
rect 15722 8146 15734 8214
rect 15484 8140 15734 8146
rect 16138 8072 17868 8430
rect 3968 6528 5088 7448
rect 3972 6322 4488 6528
rect 3034 5752 4486 6322
rect 7682 6080 7818 8050
rect 12028 6586 12928 7492
rect 6066 5984 6076 6080
rect 6770 5984 6780 6080
rect 8770 5984 8780 6080
rect 9474 5984 9484 6080
rect 3972 5544 4488 5752
rect 3972 4968 5074 5544
rect 3990 4624 5074 4968
rect 7686 4018 7818 5978
rect 12028 5488 12544 6586
rect 15544 6182 15668 7932
rect 13920 5954 13930 6050
rect 14624 5954 14634 6050
rect 16616 5960 16626 6056
rect 17320 5960 17330 6056
rect 12028 4582 12928 5488
rect 6884 3974 7514 4004
rect 6884 3722 7518 3974
rect 9376 3722 10206 3974
rect 6872 3680 10206 3722
rect 6872 3488 9804 3680
rect 10124 3564 10206 3680
rect 10124 3488 10204 3564
rect 6872 3478 10204 3488
rect 12028 3088 12544 4582
rect 15550 4124 15674 5874
rect 14466 3576 15296 3946
rect 17228 3576 18058 3936
rect 14466 3558 18452 3576
rect 18778 3558 19324 8430
rect 19874 6428 20500 9356
rect 21680 6806 22162 7214
rect 21680 6746 21738 6806
rect 21854 6746 22162 6806
rect 21680 6670 22162 6746
rect 19886 6218 20500 6428
rect 21678 6610 22162 6670
rect 21678 6556 22160 6610
rect 21678 6354 21688 6556
rect 22156 6354 22166 6556
rect 19884 6154 20502 6218
rect 19884 5792 22950 6154
rect 19884 5704 20502 5792
rect 13474 3216 13484 3470
rect 13922 3216 13932 3470
rect 12030 2956 12544 3088
rect 3020 2954 11670 2956
rect 12030 2954 12548 2956
rect 3020 2630 12548 2954
rect 13480 2876 13926 3216
rect 14466 3144 19324 3558
rect 14486 3134 19324 3144
rect 19886 2976 20500 5704
rect 20852 5206 20862 5620
rect 21408 5206 21418 5620
rect 21656 5274 21666 5674
rect 22184 5274 22194 5674
rect 20864 3242 21400 5206
rect 21052 3234 21202 3242
rect 19098 2968 20500 2976
rect 18600 2964 20506 2968
rect 14352 2916 16978 2920
rect 14352 2846 17136 2916
rect 17662 2880 20506 2964
rect 14178 2672 17136 2846
rect 3020 2394 11652 2630
rect 13490 2266 13924 2624
rect 14352 2544 17136 2672
rect 13966 2538 14114 2544
rect 13966 2496 13978 2538
rect 14102 2496 14114 2538
rect 13966 2490 14114 2496
rect 6582 2246 6754 2266
rect 6054 2240 6754 2246
rect 6054 1832 6066 2240
rect 13490 2214 13920 2266
rect 6754 1832 6756 2196
rect 13482 2162 13920 2214
rect 13482 2044 13924 2162
rect 12810 2042 13924 2044
rect 12136 1832 13924 2042
rect 6054 1824 6756 1832
rect 9598 1824 13924 1832
rect 6054 1796 13924 1824
rect 6054 1628 12994 1796
rect 6058 1522 12994 1628
rect 13490 1532 13924 1796
rect 13978 1678 14100 2490
rect 16730 2478 17136 2544
rect 17652 2742 20506 2880
rect 17652 2498 18024 2742
rect 18600 2670 20506 2742
rect 21054 2678 21192 3234
rect 21706 2850 22158 5274
rect 21706 2806 22096 2850
rect 21722 2802 21928 2806
rect 21722 2732 21734 2802
rect 21818 2732 21928 2802
rect 21722 2726 21830 2732
rect 18510 2480 19776 2516
rect 16730 2276 17406 2478
rect 18510 2442 19424 2480
rect 18298 2306 19424 2442
rect 13958 1672 14100 1678
rect 13958 1620 13970 1672
rect 14066 1622 14100 1672
rect 17646 2002 18032 2252
rect 18510 2242 19424 2306
rect 19790 2242 19800 2480
rect 21380 2378 21784 2552
rect 18510 2222 19776 2242
rect 17646 1862 17722 2002
rect 18010 1862 18032 2002
rect 17646 1714 18032 1862
rect 18098 2170 18226 2176
rect 18098 2102 18110 2170
rect 18214 2102 18226 2170
rect 18098 2096 18226 2102
rect 14066 1620 14078 1622
rect 13958 1614 14078 1620
rect 9918 1520 12994 1522
rect 9918 1516 10410 1520
rect 10646 1512 12994 1520
rect 12136 1508 12994 1512
rect 14324 1468 17306 1598
rect 17646 1542 18030 1714
rect 18098 1700 18220 2096
rect 18094 1694 18224 1700
rect 18094 1634 18106 1694
rect 18212 1634 18224 1694
rect 18094 1628 18224 1634
rect 18398 1488 20892 1698
rect 18190 1486 21138 1488
rect 18190 1484 21330 1486
rect 21384 1484 21528 2378
rect 14048 1356 17530 1468
rect 18190 1366 21528 1484
rect 18190 1360 21480 1366
rect 10878 1192 10888 1198
rect 10874 844 10888 1192
rect 11288 844 11298 1198
rect 13500 1182 13920 1262
rect 14324 1224 17306 1356
rect 18190 1352 21330 1360
rect 13500 1126 13568 1182
rect 13814 1126 13920 1182
rect 13500 970 13920 1126
rect 10874 722 11256 844
rect 13496 722 13920 970
rect 17650 1214 18048 1298
rect 18398 1234 20892 1352
rect 17650 1146 17752 1214
rect 17938 1146 18048 1214
rect 17650 1000 18048 1146
rect 21718 1130 21830 1492
rect 21702 1124 21842 1130
rect 21048 1116 21186 1122
rect 21048 1042 21060 1116
rect 21174 1042 21186 1116
rect 21702 1050 21714 1124
rect 21830 1050 21842 1124
rect 21702 1044 21842 1050
rect 21048 1036 21186 1042
rect 17650 722 18050 1000
rect 21060 970 21174 1036
rect 21718 970 21830 1044
rect 20818 722 22096 970
rect 2996 712 22096 722
rect 2996 210 22976 712
rect 2996 206 20672 210
<< via1 >>
rect 5946 11698 7362 12068
rect 5246 11342 5628 11454
rect 6478 11102 6860 11214
rect 5238 10850 5636 10954
rect 6482 10596 6864 10708
rect 5234 10334 5636 10424
rect 6488 10080 6870 10192
rect 7640 11354 8022 11466
rect 16012 11346 16350 11572
rect 8814 11088 9196 11200
rect 7640 10840 8022 10952
rect 8814 10580 9196 10692
rect 7640 10328 8022 10440
rect 8814 10066 9196 10178
rect 5226 9828 5636 9894
rect 7640 9814 8022 9926
rect 12212 10024 12602 10350
rect 7550 9306 8068 9526
rect 11414 9290 11702 9704
rect 16012 9496 16354 9736
rect 21752 10002 21852 10288
rect 21034 9684 21190 9854
rect 10382 8626 10854 8984
rect 6076 5984 6770 6080
rect 8780 5984 9474 6080
rect 13930 5954 14624 6050
rect 16626 5960 17320 6056
rect 9804 3488 10124 3680
rect 21688 6354 22156 6556
rect 13484 3216 13922 3470
rect 20862 5206 21408 5620
rect 21666 5274 22184 5674
rect 6066 1832 6754 2240
rect 19424 2242 19790 2480
rect 17722 1862 18010 2002
rect 10888 844 11288 1198
<< metal2 >>
rect 5946 12068 7362 12078
rect 5250 11938 5630 11946
rect 5676 11938 5946 11956
rect 5250 11704 5946 11938
rect 5250 11696 5862 11704
rect 7362 11938 7662 11946
rect 7362 11698 8036 11938
rect 5946 11696 8036 11698
rect 5250 11464 5630 11696
rect 5946 11694 8024 11696
rect 5946 11688 7362 11694
rect 5246 11454 5630 11464
rect 5628 11446 5630 11454
rect 7626 11466 8024 11694
rect 16012 11572 16350 11582
rect 5628 11342 5636 11446
rect 5246 11332 5636 11342
rect 5254 10964 5636 11332
rect 7626 11354 7640 11466
rect 8022 11354 8028 11466
rect 6478 11214 6860 11224
rect 5238 10954 5636 10964
rect 5238 10840 5636 10850
rect 5242 10434 5636 10840
rect 5234 10424 5636 10434
rect 5226 10334 5234 10404
rect 6472 11102 6478 11214
rect 6860 11102 6872 11214
rect 7626 11134 8028 11354
rect 16350 11346 16354 11560
rect 6472 10708 6872 11102
rect 6472 10596 6482 10708
rect 6864 10596 6872 10708
rect 6472 10338 6872 10596
rect 7632 10952 8028 11134
rect 7632 10840 7640 10952
rect 8022 10840 8028 10952
rect 7632 10440 8028 10840
rect 5226 10324 5636 10334
rect 5226 9904 5614 10324
rect 6470 10192 6878 10338
rect 6470 10080 6488 10192
rect 6870 10080 6878 10192
rect 5226 9894 5636 9904
rect 5226 9818 5636 9828
rect 6470 9526 6878 10080
rect 7632 10328 7640 10440
rect 8022 10328 8028 10440
rect 7632 9926 8028 10328
rect 7632 9814 7640 9926
rect 8022 9814 8028 9926
rect 8814 11200 9196 11210
rect 9196 11088 9206 11198
rect 8814 10692 9206 11088
rect 9196 10580 9206 10692
rect 8814 10178 9206 10580
rect 9196 10066 9206 10178
rect 7640 9804 8022 9814
rect 7550 9526 8068 9536
rect 8814 9526 9206 10066
rect 12072 10360 12472 10366
rect 12072 10350 12602 10360
rect 12072 10024 12212 10350
rect 12072 10014 12602 10024
rect 11414 9704 11702 9714
rect 6468 9306 7550 9526
rect 8068 9306 9212 9526
rect 6468 9304 9212 9306
rect 7550 9296 8068 9304
rect 11414 9280 11702 9290
rect 10382 8984 10854 8994
rect 10382 8616 10854 8626
rect 6076 6080 6770 6090
rect 8780 6086 9474 6090
rect 6070 5984 6076 6036
rect 6070 5974 6770 5984
rect 8762 6080 9488 6086
rect 8762 5984 8780 6080
rect 9474 5984 9488 6080
rect 6070 5660 6762 5974
rect 6050 5432 6768 5660
rect 6050 5404 6854 5432
rect 8762 5404 9488 5984
rect 6050 5124 9488 5404
rect 6050 5096 6854 5124
rect 6050 2240 6768 5096
rect 12072 4514 12472 10014
rect 16012 9736 16354 11346
rect 21752 10288 21852 10298
rect 19412 10018 21752 10264
rect 19412 10012 20960 10018
rect 16012 9486 16354 9496
rect 13930 6050 14624 6060
rect 13924 5954 13930 6040
rect 16626 6056 17320 6066
rect 14624 5954 14636 6040
rect 13924 5416 14636 5954
rect 16604 5960 16626 6022
rect 17320 5960 17330 6022
rect 16604 5416 17330 5960
rect 13924 5162 17330 5416
rect 13924 5152 15956 5162
rect 16174 5152 17330 5162
rect 13924 5146 14636 5152
rect 10900 4110 12472 4514
rect 10900 4108 12468 4110
rect 10900 3960 11256 4108
rect 9804 3680 10124 3690
rect 9804 3478 10124 3488
rect 6050 1998 6066 2240
rect 6754 1998 6768 2240
rect 6066 1822 6754 1832
rect 10898 1202 11258 3960
rect 13464 3490 13944 3500
rect 13464 3184 13944 3194
rect 16174 2274 16606 5152
rect 19420 2490 19784 10012
rect 21752 9992 21852 10002
rect 21034 9860 21190 9864
rect 20872 9854 21416 9860
rect 20872 9684 21034 9854
rect 21190 9684 21416 9854
rect 20872 5732 21416 9684
rect 21688 6556 22156 6566
rect 21688 5906 22156 6354
rect 20872 5630 21408 5732
rect 21688 5684 22160 5906
rect 20862 5620 21408 5630
rect 21666 5674 22184 5684
rect 21666 5264 22184 5274
rect 20862 5196 21408 5206
rect 19420 2480 19790 2490
rect 16174 2148 16604 2274
rect 19420 2256 19424 2480
rect 19424 2232 19790 2242
rect 16170 2020 17090 2148
rect 16170 2002 18038 2020
rect 16170 1862 17722 2002
rect 18010 1862 18038 2002
rect 16170 1828 18038 1862
rect 16170 1764 17090 1828
rect 10898 1198 11304 1202
rect 10838 844 10888 1198
rect 11288 1090 11304 1198
rect 10838 834 11288 844
rect 10838 826 11282 834
<< via2 >>
rect 11414 9290 11702 9704
rect 10382 8626 10854 8984
rect 9804 3488 10124 3680
rect 13464 3470 13944 3490
rect 13464 3216 13484 3470
rect 13484 3216 13922 3470
rect 13922 3216 13944 3470
rect 13464 3194 13944 3216
<< metal3 >>
rect 11404 9704 11712 9709
rect 11404 9290 11414 9704
rect 11702 9362 11712 9704
rect 11702 9290 11834 9362
rect 11404 9285 11834 9290
rect 11448 9284 11834 9285
rect 11448 9176 11835 9284
rect 10330 8990 11190 9142
rect 10330 8984 11224 8990
rect 10330 8626 10382 8984
rect 10854 8626 11224 8984
rect 10330 8348 11190 8626
rect 10878 3724 11089 8348
rect 10696 3688 11089 3724
rect 9970 3685 11089 3688
rect 9794 3680 11089 3685
rect 9794 3488 9804 3680
rect 10124 3511 11089 3680
rect 10124 3488 10912 3511
rect 11540 3490 11835 9176
rect 13454 3490 13954 3495
rect 9794 3486 10912 3488
rect 9794 3484 10572 3486
rect 11534 3484 11998 3490
rect 13454 3484 13464 3490
rect 9794 3483 10536 3484
rect 9908 3474 10536 3483
rect 11534 3194 13464 3484
rect 13944 3194 13954 3490
rect 11534 3184 11998 3194
rect 13454 3189 13954 3194
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM1
timestamp 1752660100
transform 0 1 7751 -1 0 6037
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM2
timestamp 1752660100
transform 0 1 15607 -1 0 6011
box -2225 -2837 2225 2837
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM3
timestamp 1752660100
transform 0 1 17848 -1 0 2372
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM4
timestamp 1752660100
transform 0 1 17860 -1 0 1422
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM5
timestamp 1752660100
transform 0 1 13722 -1 0 1400
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM6
timestamp 1752660100
transform 0 1 13736 -1 0 2758
box -296 -610 296 610
use sky130_fd_pr__pfet_01v8_lvt_CYPNY8  XM7
timestamp 1752660100
transform 0 1 15237 -1 0 10275
box -419 -519 419 519
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM8
timestamp 1752660100
transform 0 1 17111 -1 0 11437
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM9
timestamp 1752660100
transform 0 1 15243 -1 0 11445
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_CYPNY8  XM10
timestamp 1752660100
transform 0 1 17109 -1 0 10271
box -419 -519 419 519
use sky130_fd_pr__pfet_01v8_lvt_6VJTDW  XM11
timestamp 1752660100
transform 0 1 7282 -1 0 10644
box -936 -2332 946 2342
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR1
timestamp 1752660100
transform -1 0 21119 0 -1 2118
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1752660100
transform 0 1 11116 -1 0 11645
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR3
timestamp 1752660100
transform 0 1 11928 -1 0 10945
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_DBPYMX  XR4
timestamp 1752660100
transform -1 0 21771 0 -1 1925
box -201 -889 201 889
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR5
timestamp 1752660100
transform 1 0 22301 0 1 10878
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_Z767S8  XR6
timestamp 1752660100
transform 1 0 21797 0 1 8628
box -201 -1902 201 1902
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR7
timestamp 1752660100
transform 0 1 20436 -1 0 11485
box -201 -1082 201 1082
use sky130_fd_pr__res_xhigh_po_0p35_MAXMKG  XR8
timestamp 1752660100
transform 0 1 20136 -1 0 10707
box -201 -742 201 742
<< labels >>
flabel metal1 3278 12260 3478 12460 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 3276 426 3476 626 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 22624 5878 22824 6078 0 FreeSans 256 0 0 0 OUT
port 2 nsew
rlabel metal1 8266 8090 9996 8998 1 S
rlabel metal2 16012 9736 16354 11346 1 G
rlabel metal1 15016 10684 15466 11196 1 D9
rlabel metal1 16932 10678 17318 11188 1 D10
rlabel metal1 15598 10118 16754 10436 1 Vc2
rlabel metal1 14048 1356 17530 1468 1 Vc
rlabel metal1 14352 2544 16978 2920 1 Vc1
rlabel space 13490 1532 13924 2624 1 D1
rlabel metal1 17646 2002 18032 2252 1 D2
rlabel metal1 9722 11138 9872 11350 1 Vb
flabel metal1 3196 5942 3396 6142 0 FreeSans 480 0 0 0 INp
port 4 nsew
flabel metal1 3274 2532 3474 2732 0 FreeSans 256 0 0 0 INm
port 3 nsew
<< end >>
