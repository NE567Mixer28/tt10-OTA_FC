magic
tech sky130A
magscale 1 2
timestamp 1768581666
<< viali >>
rect 6566 11274 6804 11392
rect 10868 11272 11104 11338
rect 3892 11040 4288 11120
rect 6592 10066 6822 10136
rect 10824 10024 11098 10098
rect 1436 8166 1990 8226
rect 9338 8154 9814 8238
rect 13108 2004 13312 2084
rect 860 1438 932 1614
rect 13152 1272 13332 1340
rect 13492 754 13740 852
rect 1378 -226 1574 -136
<< metal1 >>
rect -824 12436 862 12442
rect -890 12408 862 12436
rect -890 12404 14056 12408
rect -890 11924 15456 12404
rect -890 11638 1686 11924
rect 1676 11424 1686 11638
rect 3352 11638 15456 11924
rect 3352 11424 3362 11638
rect 3884 11126 4300 11638
rect 6460 11392 6950 11638
rect 6460 11274 6566 11392
rect 6804 11274 6950 11392
rect 6460 11196 6950 11274
rect 10764 11338 11202 11638
rect 13514 11630 15456 11638
rect 10764 11272 10868 11338
rect 11104 11272 11202 11338
rect 10764 11186 11202 11272
rect 3880 11120 4300 11126
rect 3880 11040 3892 11120
rect 4288 11040 4300 11120
rect 3880 11034 4300 11040
rect 7140 11036 10538 11088
rect 1660 10928 1670 11016
rect 2120 10928 2130 11016
rect 2908 10908 2918 10984
rect 3352 10908 3362 10984
rect -238 10100 330 10868
rect 476 10650 486 10750
rect 914 10650 924 10750
rect 1668 10402 1678 10480
rect 2118 10402 2128 10480
rect 470 10148 480 10248
rect 908 10148 918 10248
rect -896 9686 330 10100
rect 1664 9862 1674 9962
rect 2110 9862 2120 9962
rect -238 9522 330 9686
rect 472 9624 482 9724
rect 910 9624 920 9724
rect 2448 9478 2578 10904
rect 7140 10826 8590 11036
rect 8994 10826 10538 11036
rect 7140 10792 10538 10826
rect 3996 10630 4006 10736
rect 4426 10630 4436 10736
rect 2908 10412 2918 10492
rect 3348 10412 3358 10492
rect 3996 10138 4006 10244
rect 4426 10138 4436 10244
rect 6490 10136 6928 10686
rect 6490 10066 6592 10136
rect 6822 10066 6928 10136
rect 6490 9974 6928 10066
rect 10670 10098 11240 10694
rect 10670 10024 10824 10098
rect 11098 10024 11240 10098
rect 2920 9890 2930 9970
rect 3360 9890 3370 9970
rect 10670 9952 11240 10024
rect 15016 9998 15440 10014
rect 4000 9606 4010 9712
rect 4430 9606 4440 9712
rect 7202 9546 10522 9878
rect 11448 9518 15440 9998
rect 11448 9512 15230 9518
rect 1668 9374 1678 9448
rect 2106 9374 2116 9448
rect 2918 9372 2928 9452
rect 3358 9372 3368 9452
rect 6526 9442 6536 9512
rect 7006 9442 7016 9512
rect 10686 9448 11216 9456
rect 10686 9246 11290 9448
rect 13920 9246 14286 9284
rect 10686 9006 14286 9246
rect 10688 8950 14286 9006
rect 1426 8232 1436 8262
rect 1424 8160 1436 8232
rect 1426 8140 1436 8160
rect 2004 8140 2014 8262
rect 9326 8238 9826 8244
rect 9326 8154 9338 8238
rect 9814 8154 9826 8238
rect 9326 8148 9826 8154
rect 620 7996 630 8124
rect 932 7996 942 8124
rect 1274 8036 1284 8108
rect 2162 8036 2172 8108
rect 3332 8004 3342 8130
rect 3698 8004 3708 8130
rect 3990 8020 4000 8132
rect 4838 8020 4848 8132
rect 8478 8012 8488 8120
rect 8810 8012 8820 8120
rect 9094 8022 9104 8120
rect 10242 8022 10252 8120
rect 11276 8016 11286 8124
rect 11608 8016 11618 8124
rect 11834 8038 11844 8136
rect 12982 8038 12992 8136
rect -456 7730 -48 7736
rect -456 6438 332 7730
rect -456 6322 -48 6438
rect 2962 6432 3066 7726
rect -898 5800 -48 6322
rect 7464 6218 8260 7818
rect 10868 6226 10990 7832
rect 13920 6996 14286 8950
rect 13920 6644 14290 6996
rect 1156 5892 1166 6088
rect 1582 5892 1592 6088
rect 4292 5938 4302 6072
rect 4812 5938 4822 6072
rect -466 5714 -48 5800
rect 7464 5828 7930 6218
rect 10098 5896 10108 6076
rect 10564 5896 10574 6076
rect 11864 5894 11874 6062
rect 12420 5894 12430 6062
rect -466 4276 344 5714
rect -404 4266 344 4276
rect 2960 4268 3078 5714
rect 7464 4194 8274 5828
rect 10888 4222 10970 5842
rect 13924 5666 14290 6644
rect 13924 5284 15430 5666
rect 630 3922 640 4020
rect 928 3922 938 4020
rect 3324 3906 3334 4032
rect 3690 3906 3700 4032
rect -724 3380 6056 3384
rect -898 3378 6056 3380
rect 7464 3378 7930 4194
rect 8450 3918 8460 4026
rect 8782 3918 8792 4026
rect 11288 3918 11298 4026
rect 11620 3918 11630 4026
rect 13924 3522 14290 5284
rect 13924 3510 14096 3522
rect -898 2784 7930 3378
rect -724 2780 7930 2784
rect 5754 2774 7930 2780
rect 13372 3236 14096 3510
rect 14390 3236 14400 3522
rect 13372 3184 14290 3236
rect 13372 3182 14282 3184
rect 13372 2392 13806 3182
rect 11660 2358 11966 2376
rect 11660 2220 13130 2358
rect 11660 1704 11966 2220
rect 13446 2114 13456 2198
rect 13726 2114 13736 2198
rect 14024 2136 15376 2468
rect 13096 2084 13324 2090
rect 13096 2004 13108 2084
rect 13312 2004 13324 2084
rect 13096 1998 13324 2004
rect 1294 1630 1304 1696
rect 1650 1630 1660 1696
rect 854 1614 938 1626
rect 854 1590 860 1614
rect 588 1440 860 1590
rect -64 592 -54 842
rect 388 592 398 842
rect 588 -352 790 1440
rect 854 1438 860 1440
rect 932 1438 938 1614
rect 2202 1610 11970 1704
rect 1898 1462 11970 1610
rect 854 1426 938 1438
rect 1276 1370 1286 1432
rect 1676 1370 1686 1432
rect 2202 1306 11970 1462
rect 13114 1346 13324 1998
rect 13114 1340 13344 1346
rect 13114 1276 13152 1340
rect 13140 1272 13152 1276
rect 13332 1272 13344 1340
rect 13140 1266 13344 1272
rect 13930 1238 15282 1240
rect 13476 1152 13486 1232
rect 13732 1152 13742 1232
rect 12458 998 13262 1104
rect 1266 162 1276 224
rect 1666 162 1676 224
rect 1814 112 2396 116
rect 1814 -26 2400 112
rect 1274 -136 1682 -58
rect 1274 -226 1378 -136
rect 1574 -226 1682 -136
rect 1274 -352 1682 -226
rect 588 -516 1682 -352
rect 738 -518 1682 -516
rect 1274 -2724 1682 -518
rect 2132 -378 2400 -26
rect 12458 -378 12806 998
rect 13436 852 13758 948
rect 13930 908 15376 1238
rect 15028 904 15376 908
rect 13436 754 13492 852
rect 13740 754 13758 852
rect 2132 -792 12808 -378
rect 2132 -802 2400 -792
rect 13436 -2724 13758 754
rect 592 -2730 14028 -2724
rect -914 -2732 14028 -2730
rect -914 -2860 15444 -2732
rect -908 -3494 15444 -2860
rect -908 -3496 972 -3494
rect -908 -3502 -536 -3496
<< via1 >>
rect 1686 11424 3352 11924
rect 1670 10928 2120 11016
rect 2918 10908 3352 10984
rect 486 10650 914 10750
rect 1678 10402 2118 10480
rect 480 10148 908 10248
rect 1674 9862 2110 9962
rect 482 9624 910 9724
rect 8590 10826 8994 11036
rect 4006 10630 4426 10736
rect 2918 10412 3348 10492
rect 4006 10138 4426 10244
rect 2930 9890 3360 9970
rect 4010 9606 4430 9712
rect 1678 9374 2106 9448
rect 2928 9372 3358 9452
rect 6536 9442 7006 9512
rect 1436 8226 2004 8262
rect 1436 8166 1990 8226
rect 1990 8166 2004 8226
rect 1436 8140 2004 8166
rect 9338 8154 9814 8238
rect 630 7996 932 8124
rect 1284 8036 2162 8108
rect 3342 8004 3698 8130
rect 4000 8020 4838 8132
rect 8488 8012 8810 8120
rect 9104 8022 10242 8120
rect 11286 8016 11608 8124
rect 11844 8038 12982 8136
rect 1166 5892 1582 6088
rect 4302 5938 4812 6072
rect 10108 5896 10564 6076
rect 11874 5894 12420 6062
rect 640 3922 928 4020
rect 3334 3906 3690 4032
rect 8460 3918 8782 4026
rect 11298 3918 11620 4026
rect 14096 3236 14390 3522
rect 13456 2114 13726 2198
rect 1304 1630 1650 1696
rect -54 592 388 842
rect 1286 1370 1676 1432
rect 13486 1152 13732 1232
rect 1276 162 1666 224
<< metal2 >>
rect 1686 11924 3352 11934
rect 1686 11414 3352 11424
rect 1688 11026 2106 11414
rect 1670 11016 2120 11026
rect 2930 10994 3352 11414
rect 1670 10918 2120 10928
rect 2918 10984 3352 10994
rect 486 10750 918 10798
rect 914 10650 918 10750
rect 486 10258 918 10650
rect 480 10248 918 10258
rect 908 10148 918 10248
rect 480 10138 918 10148
rect 486 9734 918 10138
rect 482 9724 918 9734
rect 910 9624 918 9724
rect 482 9614 918 9624
rect 486 9136 918 9614
rect 1674 10490 2114 10918
rect 2918 10898 3352 10908
rect 2930 10502 3352 10898
rect 8590 11036 8994 11046
rect 8590 10816 8994 10826
rect 4006 10736 4426 10746
rect 4006 10620 4426 10630
rect 2918 10492 3352 10502
rect 1674 10480 2118 10490
rect 1674 10402 1678 10480
rect 3348 10412 3352 10492
rect 2918 10402 3352 10412
rect 1674 10392 2118 10402
rect 1674 9962 2114 10392
rect 2110 9862 2114 9962
rect 1674 9448 2114 9862
rect 2930 9980 3352 10402
rect 4012 10254 4412 10620
rect 4006 10244 4426 10254
rect 4006 10128 4426 10138
rect 2930 9970 3360 9980
rect 2930 9880 3360 9890
rect 2930 9462 3352 9880
rect 4012 9722 4412 10128
rect 4010 9712 4430 9722
rect 4010 9596 4430 9606
rect 1674 9374 1678 9448
rect 2106 9374 2114 9448
rect 1674 9356 2114 9374
rect 2928 9452 3358 9462
rect 2928 9362 3358 9372
rect 2930 9352 3352 9362
rect 4012 9136 4412 9596
rect 6536 9512 7006 9522
rect 6536 9432 7006 9442
rect 486 9002 4412 9136
rect 494 8840 4412 9002
rect 494 8784 12718 8840
rect 494 8736 13030 8784
rect 1136 8262 2290 8736
rect 1136 8140 1436 8262
rect 2004 8140 2290 8262
rect 3852 8462 13030 8736
rect 630 8124 932 8134
rect 1136 8108 2290 8140
rect 1136 8072 1284 8108
rect 2162 8072 2290 8108
rect 3342 8130 3698 8140
rect 1284 8026 2162 8036
rect 630 7986 932 7996
rect 3852 8132 5006 8462
rect 3852 8064 4000 8132
rect 4838 8064 5006 8132
rect 8964 8238 10306 8462
rect 8964 8154 9338 8238
rect 9814 8154 10306 8238
rect 8488 8120 8810 8130
rect 4000 8010 4838 8020
rect 8472 8012 8488 8120
rect 8964 8120 10306 8154
rect 11688 8136 13030 8462
rect 8964 8052 9104 8120
rect 10242 8052 10306 8120
rect 11286 8124 11608 8134
rect 9104 8012 10242 8022
rect 11268 8016 11286 8104
rect 11688 8044 11844 8136
rect 12982 8044 13030 8136
rect 11844 8028 12982 8038
rect 3342 7994 3698 8004
rect 8472 8002 8810 8012
rect 11268 8006 11608 8016
rect 652 4030 916 7986
rect 1166 6088 1582 6098
rect 640 4020 928 4030
rect 640 3912 928 3922
rect 1166 3332 1582 5892
rect 3352 4042 3658 7994
rect 4302 6072 4812 6082
rect 4302 5928 4812 5938
rect 3334 4032 3690 4042
rect 3334 3896 3690 3906
rect 4338 3332 4774 5928
rect 8472 4036 8806 8002
rect 10108 6076 10564 6086
rect 10564 5896 10594 6024
rect 10108 5886 10594 5896
rect 8460 4026 8806 4036
rect 8782 3930 8806 4026
rect 8460 3908 8782 3918
rect 10138 3622 10594 5886
rect 11268 4036 11602 8006
rect 11874 6062 12420 6072
rect 11874 5884 12420 5894
rect 11268 4026 11620 4036
rect 11268 3918 11298 4026
rect 11268 3914 11620 3918
rect 11298 3908 11620 3914
rect 11894 3640 12366 5884
rect 11894 3622 12752 3640
rect 10138 3382 12752 3622
rect 1166 2912 4774 3332
rect 10152 3254 12752 3382
rect 12226 3248 12752 3254
rect 1166 2904 4752 2912
rect 1166 2594 1582 2904
rect -586 2336 1582 2594
rect -586 2162 1578 2336
rect -586 1158 -58 2162
rect 12250 1912 12752 3248
rect 14096 3522 14390 3532
rect 14096 3226 14390 3236
rect 13456 2198 13726 2208
rect 13368 2114 13456 2180
rect 13726 2114 13818 2180
rect 13368 1912 13818 2114
rect 1304 1696 1650 1706
rect 1304 1620 1650 1630
rect 12250 1516 13878 1912
rect 12562 1508 13878 1516
rect 1286 1432 1676 1442
rect 1266 1370 1286 1412
rect 1266 1360 1676 1370
rect 1266 1158 1668 1360
rect 13368 1232 13818 1508
rect 13368 1182 13486 1232
rect -586 842 1734 1158
rect 13732 1182 13818 1232
rect 13486 1142 13732 1152
rect -586 592 -54 842
rect 388 592 1734 842
rect -586 542 1734 592
rect -572 534 1734 542
rect 1266 224 1668 534
rect 1266 178 1276 224
rect 1666 178 1668 224
rect 1276 152 1666 162
<< via2 >>
rect 8590 10826 8994 11036
rect 6536 9442 7006 9512
rect 14096 3236 14390 3522
rect 1304 1630 1650 1696
rect -54 592 388 842
<< metal3 >>
rect 8580 11036 9004 11041
rect 8580 10826 8590 11036
rect 8994 10826 9004 11036
rect 8580 10821 9004 10826
rect 6526 9512 7016 9517
rect 6526 9486 6536 9512
rect 6442 9442 6536 9486
rect 7006 9486 7016 9512
rect 7006 9442 7054 9486
rect 6442 9216 7054 9442
rect 8616 9216 8954 10821
rect 6442 9188 8954 9216
rect 6436 9038 8954 9188
rect 6436 9000 7054 9038
rect 8616 9030 8954 9038
rect 1310 3282 1896 3292
rect 6436 3282 7038 9000
rect 1310 2896 7038 3282
rect 14086 3522 14400 3527
rect 14086 3236 14096 3522
rect 14390 3236 14400 3522
rect 14086 3231 14400 3236
rect 1310 2884 6754 2896
rect 1310 1701 1896 2884
rect 1294 1696 1896 1701
rect 1294 1630 1304 1696
rect 1650 1646 1896 1696
rect 1650 1630 1660 1646
rect 1294 1625 1660 1630
rect -64 842 398 847
rect -64 592 -54 842
rect 388 592 398 842
rect -64 587 398 592
<< via3 >>
rect 14096 3236 14390 3522
rect -54 592 388 842
<< metal4 >>
rect 14182 3556 14552 3560
rect 14182 3523 14730 3556
rect 14095 3522 14730 3523
rect 14095 3236 14096 3522
rect 14390 3236 14730 3522
rect 14095 3235 14730 3236
rect 14182 3180 14730 3235
rect -55 842 389 843
rect -55 592 -54 842
rect 388 592 389 842
rect -55 591 389 592
rect -22 -2030 328 591
rect 14356 478 14730 3180
rect 13988 468 14730 478
rect 12022 466 14730 468
rect 11844 170 14730 466
rect 11844 166 12156 170
rect 13988 166 14730 170
rect 798 -2030 2386 -2018
rect -22 -2430 2386 -2030
rect -22 -2442 328 -2430
use sky130_fd_pr__cap_mim_m3_1_7MGYMT  XC1
timestamp 1768572465
transform 0 1 7104 -1 0 152
box -2426 -4800 2426 4800
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM1
timestamp 1768572465
transform 0 1 3019 -1 0 6019
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_lvt_BFTKM6  XM2
timestamp 1768572465
transform 0 1 10939 -1 0 6019
box -2225 -2837 2225 2837
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM3
timestamp 1768572465
transform 0 1 13576 -1 0 2288
box -296 -610 296 610
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM4
timestamp 1768572465
transform 0 1 13600 -1 0 1056
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_WVASGV  XM5
timestamp 1768572465
transform 0 1 1474 -1 0 64
box -296 -490 296 490
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM6
timestamp 1768572465
transform 0 1 1452 -1 0 1534
box -296 -610 296 610
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM7
timestamp 1768572465
transform 0 1 6731 -1 0 9733
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_EABQL5  XM8
timestamp 1768572465
transform 0 1 10978 -1 0 10939
box -419 -604 419 604
use sky130_fd_pr__pfet_01v8_lvt_EABQL5  XM9
timestamp 1768572465
transform 0 1 6706 -1 0 10949
box -419 -604 419 604
use sky130_fd_pr__pfet_01v8_lvt_2L7S3R  XM10
timestamp 1768572465
transform 0 1 10971 -1 0 9701
box -419 -619 419 619
use sky130_fd_pr__pfet_01v8_lvt_6VJTDW  XM11
timestamp 1768572465
transform 0 1 2513 -1 0 10189
box -941 -2337 941 2337
<< labels >>
flabel metal1 -846 5978 -646 6178 0 FreeSans 256 0 0 0 INp
port 5 nsew
flabel metal1 -846 3022 -646 3222 0 FreeSans 256 0 0 0 INm
port 6 nsew
flabel metal1 -856 9790 -656 9990 0 FreeSans 256 0 0 0 Vb
port 0 nsew
flabel metal1 15156 5378 15356 5578 0 FreeSans 256 0 0 0 OUT
port 4 nsew
flabel metal1 15156 2190 15356 2390 0 FreeSans 256 0 0 0 Vc1
port 7 nsew
flabel metal1 15150 978 15350 1178 0 FreeSans 256 0 0 0 Vc
port 8 nsew
flabel metal1 15148 9736 15348 9936 0 FreeSans 256 0 0 0 Vc2
port 3 nsew
flabel metal1 -812 11902 -612 12102 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 -826 -3208 -626 -3008 0 FreeSans 256 0 0 0 GND
port 2 nsew
rlabel metal2 12250 1516 12752 3640 1 D2
rlabel metal2 -586 542 -58 2594 1 D1
rlabel metal3 8616 9030 8954 10826 1 G
rlabel metal1 6490 10136 6928 10686 1 D9
rlabel metal1 10670 10098 11240 10694 1 D10
rlabel metal2 3852 8132 5006 8840 1 S
<< end >>
